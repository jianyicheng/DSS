module STORE_QUEUE_LSQ_A( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_8, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_9, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_10, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_11, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_12, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_13, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_14, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_15, // @[:@6.4]
  input         io_bbNumStores, // @[:@6.4]
  output [3:0]  io_storeTail, // @[:@6.4]
  output [3:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [3:0]  io_loadTail, // @[:@6.4]
  input  [3:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadAddressDone_8, // @[:@6.4]
  input         io_loadAddressDone_9, // @[:@6.4]
  input         io_loadAddressDone_10, // @[:@6.4]
  input         io_loadAddressDone_11, // @[:@6.4]
  input         io_loadAddressDone_12, // @[:@6.4]
  input         io_loadAddressDone_13, // @[:@6.4]
  input         io_loadAddressDone_14, // @[:@6.4]
  input         io_loadAddressDone_15, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input         io_loadDataDone_8, // @[:@6.4]
  input         io_loadDataDone_9, // @[:@6.4]
  input         io_loadDataDone_10, // @[:@6.4]
  input         io_loadDataDone_11, // @[:@6.4]
  input         io_loadDataDone_12, // @[:@6.4]
  input         io_loadDataDone_13, // @[:@6.4]
  input         io_loadDataDone_14, // @[:@6.4]
  input         io_loadDataDone_15, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_7, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_8, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_9, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_10, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_11, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_12, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_13, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_14, // @[:@6.4]
  input  [31:0] io_loadAddressQueue_15, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeAddrDone_8, // @[:@6.4]
  output        io_storeAddrDone_9, // @[:@6.4]
  output        io_storeAddrDone_10, // @[:@6.4]
  output        io_storeAddrDone_11, // @[:@6.4]
  output        io_storeAddrDone_12, // @[:@6.4]
  output        io_storeAddrDone_13, // @[:@6.4]
  output        io_storeAddrDone_14, // @[:@6.4]
  output        io_storeAddrDone_15, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output        io_storeDataDone_8, // @[:@6.4]
  output        io_storeDataDone_9, // @[:@6.4]
  output        io_storeDataDone_10, // @[:@6.4]
  output        io_storeDataDone_11, // @[:@6.4]
  output        io_storeDataDone_12, // @[:@6.4]
  output        io_storeDataDone_13, // @[:@6.4]
  output        io_storeDataDone_14, // @[:@6.4]
  output        io_storeDataDone_15, // @[:@6.4]
  output [31:0] io_storeAddrQueue_0, // @[:@6.4]
  output [31:0] io_storeAddrQueue_1, // @[:@6.4]
  output [31:0] io_storeAddrQueue_2, // @[:@6.4]
  output [31:0] io_storeAddrQueue_3, // @[:@6.4]
  output [31:0] io_storeAddrQueue_4, // @[:@6.4]
  output [31:0] io_storeAddrQueue_5, // @[:@6.4]
  output [31:0] io_storeAddrQueue_6, // @[:@6.4]
  output [31:0] io_storeAddrQueue_7, // @[:@6.4]
  output [31:0] io_storeAddrQueue_8, // @[:@6.4]
  output [31:0] io_storeAddrQueue_9, // @[:@6.4]
  output [31:0] io_storeAddrQueue_10, // @[:@6.4]
  output [31:0] io_storeAddrQueue_11, // @[:@6.4]
  output [31:0] io_storeAddrQueue_12, // @[:@6.4]
  output [31:0] io_storeAddrQueue_13, // @[:@6.4]
  output [31:0] io_storeAddrQueue_14, // @[:@6.4]
  output [31:0] io_storeAddrQueue_15, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_8, // @[:@6.4]
  output [31:0] io_storeDataQueue_9, // @[:@6.4]
  output [31:0] io_storeDataQueue_10, // @[:@6.4]
  output [31:0] io_storeDataQueue_11, // @[:@6.4]
  output [31:0] io_storeDataQueue_12, // @[:@6.4]
  output [31:0] io_storeDataQueue_13, // @[:@6.4]
  output [31:0] io_storeDataQueue_14, // @[:@6.4]
  output [31:0] io_storeDataQueue_15, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input  [31:0] io_addressFromStorePorts_0, // @[:@6.4]
  output [31:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  output        io_storeEnableToMem, // @[:@6.4]
  input         io_memIsReadyForStores // @[:@6.4]
);
  reg [3:0] head; // @[StoreQueue.scala 50:21:@8.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[StoreQueue.scala 51:21:@9.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[StoreQueue.scala 53:24:@27.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[StoreQueue.scala 54:22:@45.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[StoreQueue.scala 55:22:@63.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[StoreQueue.scala 56:22:@81.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[StoreQueue.scala 57:26:@99.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[StoreQueue.scala 58:26:@117.4]
  reg [31:0] _RAND_97;
  reg  allocatedEntries_0; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_98;
  reg  allocatedEntries_1; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_99;
  reg  allocatedEntries_2; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_100;
  reg  allocatedEntries_3; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_101;
  reg  allocatedEntries_4; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_102;
  reg  allocatedEntries_5; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_103;
  reg  allocatedEntries_6; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_104;
  reg  allocatedEntries_7; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_105;
  reg  allocatedEntries_8; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_106;
  reg  allocatedEntries_9; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_107;
  reg  allocatedEntries_10; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_108;
  reg  allocatedEntries_11; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_109;
  reg  allocatedEntries_12; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_110;
  reg  allocatedEntries_13; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_111;
  reg  allocatedEntries_14; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_112;
  reg  allocatedEntries_15; // @[StoreQueue.scala 59:33:@135.4]
  reg [31:0] _RAND_113;
  reg  storeCompleted_0; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_114;
  reg  storeCompleted_1; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_115;
  reg  storeCompleted_2; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_116;
  reg  storeCompleted_3; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_117;
  reg  storeCompleted_4; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_118;
  reg  storeCompleted_5; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_119;
  reg  storeCompleted_6; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_120;
  reg  storeCompleted_7; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_121;
  reg  storeCompleted_8; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_122;
  reg  storeCompleted_9; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_123;
  reg  storeCompleted_10; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_124;
  reg  storeCompleted_11; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_125;
  reg  storeCompleted_12; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_126;
  reg  storeCompleted_13; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_127;
  reg  storeCompleted_14; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_128;
  reg  storeCompleted_15; // @[StoreQueue.scala 60:31:@153.4]
  reg [31:0] _RAND_129;
  reg  checkBits_0; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_130;
  reg  checkBits_1; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_131;
  reg  checkBits_2; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_132;
  reg  checkBits_3; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_133;
  reg  checkBits_4; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_134;
  reg  checkBits_5; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_135;
  reg  checkBits_6; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_136;
  reg  checkBits_7; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_137;
  reg  checkBits_8; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_138;
  reg  checkBits_9; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_139;
  reg  checkBits_10; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_140;
  reg  checkBits_11; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_141;
  reg  checkBits_12; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_142;
  reg  checkBits_13; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_143;
  reg  checkBits_14; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_144;
  reg  checkBits_15; // @[StoreQueue.scala 61:26:@171.4]
  reg [31:0] _RAND_145;
  wire [5:0] _GEN_1138; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1596; // @[util.scala 14:20:@173.4]
  wire [6:0] _T_1597; // @[util.scala 14:20:@174.4]
  wire [5:0] _T_1598; // @[util.scala 14:20:@175.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@176.4]
  wire [4:0] _T_1599; // @[util.scala 14:25:@176.4]
  wire [4:0] _GEN_1139; // @[StoreQueue.scala 70:46:@177.4]
  wire  _T_1600; // @[StoreQueue.scala 70:46:@177.4]
  wire  initBits_0; // @[StoreQueue.scala 70:64:@178.4]
  wire [6:0] _T_1605; // @[util.scala 14:20:@180.4]
  wire [6:0] _T_1606; // @[util.scala 14:20:@181.4]
  wire [5:0] _T_1607; // @[util.scala 14:20:@182.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@183.4]
  wire [4:0] _T_1608; // @[util.scala 14:25:@183.4]
  wire  _T_1609; // @[StoreQueue.scala 70:46:@184.4]
  wire  initBits_1; // @[StoreQueue.scala 70:64:@185.4]
  wire [6:0] _T_1614; // @[util.scala 14:20:@187.4]
  wire [6:0] _T_1615; // @[util.scala 14:20:@188.4]
  wire [5:0] _T_1616; // @[util.scala 14:20:@189.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@190.4]
  wire [4:0] _T_1617; // @[util.scala 14:25:@190.4]
  wire  _T_1618; // @[StoreQueue.scala 70:46:@191.4]
  wire  initBits_2; // @[StoreQueue.scala 70:64:@192.4]
  wire [6:0] _T_1623; // @[util.scala 14:20:@194.4]
  wire [6:0] _T_1624; // @[util.scala 14:20:@195.4]
  wire [5:0] _T_1625; // @[util.scala 14:20:@196.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@197.4]
  wire [4:0] _T_1626; // @[util.scala 14:25:@197.4]
  wire  _T_1627; // @[StoreQueue.scala 70:46:@198.4]
  wire  initBits_3; // @[StoreQueue.scala 70:64:@199.4]
  wire [6:0] _T_1632; // @[util.scala 14:20:@201.4]
  wire [6:0] _T_1633; // @[util.scala 14:20:@202.4]
  wire [5:0] _T_1634; // @[util.scala 14:20:@203.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@204.4]
  wire [4:0] _T_1635; // @[util.scala 14:25:@204.4]
  wire  _T_1636; // @[StoreQueue.scala 70:46:@205.4]
  wire  initBits_4; // @[StoreQueue.scala 70:64:@206.4]
  wire [6:0] _T_1641; // @[util.scala 14:20:@208.4]
  wire [6:0] _T_1642; // @[util.scala 14:20:@209.4]
  wire [5:0] _T_1643; // @[util.scala 14:20:@210.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@211.4]
  wire [4:0] _T_1644; // @[util.scala 14:25:@211.4]
  wire  _T_1645; // @[StoreQueue.scala 70:46:@212.4]
  wire  initBits_5; // @[StoreQueue.scala 70:64:@213.4]
  wire [6:0] _T_1650; // @[util.scala 14:20:@215.4]
  wire [6:0] _T_1651; // @[util.scala 14:20:@216.4]
  wire [5:0] _T_1652; // @[util.scala 14:20:@217.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@218.4]
  wire [4:0] _T_1653; // @[util.scala 14:25:@218.4]
  wire  _T_1654; // @[StoreQueue.scala 70:46:@219.4]
  wire  initBits_6; // @[StoreQueue.scala 70:64:@220.4]
  wire [6:0] _T_1659; // @[util.scala 14:20:@222.4]
  wire [6:0] _T_1660; // @[util.scala 14:20:@223.4]
  wire [5:0] _T_1661; // @[util.scala 14:20:@224.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@225.4]
  wire [4:0] _T_1662; // @[util.scala 14:25:@225.4]
  wire  _T_1663; // @[StoreQueue.scala 70:46:@226.4]
  wire  initBits_7; // @[StoreQueue.scala 70:64:@227.4]
  wire [6:0] _T_1668; // @[util.scala 14:20:@229.4]
  wire [6:0] _T_1669; // @[util.scala 14:20:@230.4]
  wire [5:0] _T_1670; // @[util.scala 14:20:@231.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@232.4]
  wire [4:0] _T_1671; // @[util.scala 14:25:@232.4]
  wire  _T_1672; // @[StoreQueue.scala 70:46:@233.4]
  wire  initBits_8; // @[StoreQueue.scala 70:64:@234.4]
  wire [6:0] _T_1677; // @[util.scala 14:20:@236.4]
  wire [6:0] _T_1678; // @[util.scala 14:20:@237.4]
  wire [5:0] _T_1679; // @[util.scala 14:20:@238.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@239.4]
  wire [4:0] _T_1680; // @[util.scala 14:25:@239.4]
  wire  _T_1681; // @[StoreQueue.scala 70:46:@240.4]
  wire  initBits_9; // @[StoreQueue.scala 70:64:@241.4]
  wire [6:0] _T_1686; // @[util.scala 14:20:@243.4]
  wire [6:0] _T_1687; // @[util.scala 14:20:@244.4]
  wire [5:0] _T_1688; // @[util.scala 14:20:@245.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@246.4]
  wire [4:0] _T_1689; // @[util.scala 14:25:@246.4]
  wire  _T_1690; // @[StoreQueue.scala 70:46:@247.4]
  wire  initBits_10; // @[StoreQueue.scala 70:64:@248.4]
  wire [6:0] _T_1695; // @[util.scala 14:20:@250.4]
  wire [6:0] _T_1696; // @[util.scala 14:20:@251.4]
  wire [5:0] _T_1697; // @[util.scala 14:20:@252.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@253.4]
  wire [4:0] _T_1698; // @[util.scala 14:25:@253.4]
  wire  _T_1699; // @[StoreQueue.scala 70:46:@254.4]
  wire  initBits_11; // @[StoreQueue.scala 70:64:@255.4]
  wire [6:0] _T_1704; // @[util.scala 14:20:@257.4]
  wire [6:0] _T_1705; // @[util.scala 14:20:@258.4]
  wire [5:0] _T_1706; // @[util.scala 14:20:@259.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@260.4]
  wire [4:0] _T_1707; // @[util.scala 14:25:@260.4]
  wire  _T_1708; // @[StoreQueue.scala 70:46:@261.4]
  wire  initBits_12; // @[StoreQueue.scala 70:64:@262.4]
  wire [6:0] _T_1713; // @[util.scala 14:20:@264.4]
  wire [6:0] _T_1714; // @[util.scala 14:20:@265.4]
  wire [5:0] _T_1715; // @[util.scala 14:20:@266.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@267.4]
  wire [4:0] _T_1716; // @[util.scala 14:25:@267.4]
  wire  _T_1717; // @[StoreQueue.scala 70:46:@268.4]
  wire  initBits_13; // @[StoreQueue.scala 70:64:@269.4]
  wire [6:0] _T_1722; // @[util.scala 14:20:@271.4]
  wire [6:0] _T_1723; // @[util.scala 14:20:@272.4]
  wire [5:0] _T_1724; // @[util.scala 14:20:@273.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@274.4]
  wire [4:0] _T_1725; // @[util.scala 14:25:@274.4]
  wire  _T_1726; // @[StoreQueue.scala 70:46:@275.4]
  wire  initBits_14; // @[StoreQueue.scala 70:64:@276.4]
  wire [6:0] _T_1731; // @[util.scala 14:20:@278.4]
  wire [6:0] _T_1732; // @[util.scala 14:20:@279.4]
  wire [5:0] _T_1733; // @[util.scala 14:20:@280.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@281.4]
  wire [4:0] _T_1734; // @[util.scala 14:25:@281.4]
  wire  _T_1735; // @[StoreQueue.scala 70:46:@282.4]
  wire  initBits_15; // @[StoreQueue.scala 70:64:@283.4]
  wire  _T_1758; // @[StoreQueue.scala 72:78:@301.4]
  wire  _T_1759; // @[StoreQueue.scala 72:78:@302.4]
  wire  _T_1760; // @[StoreQueue.scala 72:78:@303.4]
  wire  _T_1761; // @[StoreQueue.scala 72:78:@304.4]
  wire  _T_1762; // @[StoreQueue.scala 72:78:@305.4]
  wire  _T_1763; // @[StoreQueue.scala 72:78:@306.4]
  wire  _T_1764; // @[StoreQueue.scala 72:78:@307.4]
  wire  _T_1765; // @[StoreQueue.scala 72:78:@308.4]
  wire  _T_1766; // @[StoreQueue.scala 72:78:@309.4]
  wire  _T_1767; // @[StoreQueue.scala 72:78:@310.4]
  wire  _T_1768; // @[StoreQueue.scala 72:78:@311.4]
  wire  _T_1769; // @[StoreQueue.scala 72:78:@312.4]
  wire  _T_1770; // @[StoreQueue.scala 72:78:@313.4]
  wire  _T_1771; // @[StoreQueue.scala 72:78:@314.4]
  wire  _T_1772; // @[StoreQueue.scala 72:78:@315.4]
  wire  _T_1773; // @[StoreQueue.scala 72:78:@316.4]
  wire [3:0] _T_1804; // @[:@356.6]
  wire [3:0] _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_15; // @[StoreQueue.scala 76:20:@357.6]
  wire [3:0] _GEN_32; // @[StoreQueue.scala 75:25:@350.4]
  wire  _GEN_33; // @[StoreQueue.scala 75:25:@350.4]
  wire [3:0] _T_1822; // @[:@372.6]
  wire [3:0] _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_49; // @[StoreQueue.scala 76:20:@373.6]
  wire [3:0] _GEN_66; // @[StoreQueue.scala 75:25:@366.4]
  wire  _GEN_67; // @[StoreQueue.scala 75:25:@366.4]
  wire [3:0] _T_1840; // @[:@388.6]
  wire [3:0] _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_83; // @[StoreQueue.scala 76:20:@389.6]
  wire [3:0] _GEN_100; // @[StoreQueue.scala 75:25:@382.4]
  wire  _GEN_101; // @[StoreQueue.scala 75:25:@382.4]
  wire [3:0] _T_1858; // @[:@404.6]
  wire [3:0] _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_117; // @[StoreQueue.scala 76:20:@405.6]
  wire [3:0] _GEN_134; // @[StoreQueue.scala 75:25:@398.4]
  wire  _GEN_135; // @[StoreQueue.scala 75:25:@398.4]
  wire [3:0] _T_1876; // @[:@420.6]
  wire [3:0] _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_151; // @[StoreQueue.scala 76:20:@421.6]
  wire [3:0] _GEN_168; // @[StoreQueue.scala 75:25:@414.4]
  wire  _GEN_169; // @[StoreQueue.scala 75:25:@414.4]
  wire [3:0] _T_1894; // @[:@436.6]
  wire [3:0] _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_185; // @[StoreQueue.scala 76:20:@437.6]
  wire [3:0] _GEN_202; // @[StoreQueue.scala 75:25:@430.4]
  wire  _GEN_203; // @[StoreQueue.scala 75:25:@430.4]
  wire [3:0] _T_1912; // @[:@452.6]
  wire [3:0] _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_219; // @[StoreQueue.scala 76:20:@453.6]
  wire [3:0] _GEN_236; // @[StoreQueue.scala 75:25:@446.4]
  wire  _GEN_237; // @[StoreQueue.scala 75:25:@446.4]
  wire [3:0] _T_1930; // @[:@468.6]
  wire [3:0] _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_253; // @[StoreQueue.scala 76:20:@469.6]
  wire [3:0] _GEN_270; // @[StoreQueue.scala 75:25:@462.4]
  wire  _GEN_271; // @[StoreQueue.scala 75:25:@462.4]
  wire [3:0] _T_1948; // @[:@484.6]
  wire [3:0] _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_287; // @[StoreQueue.scala 76:20:@485.6]
  wire [3:0] _GEN_304; // @[StoreQueue.scala 75:25:@478.4]
  wire  _GEN_305; // @[StoreQueue.scala 75:25:@478.4]
  wire [3:0] _T_1966; // @[:@500.6]
  wire [3:0] _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_321; // @[StoreQueue.scala 76:20:@501.6]
  wire [3:0] _GEN_338; // @[StoreQueue.scala 75:25:@494.4]
  wire  _GEN_339; // @[StoreQueue.scala 75:25:@494.4]
  wire [3:0] _T_1984; // @[:@516.6]
  wire [3:0] _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_355; // @[StoreQueue.scala 76:20:@517.6]
  wire [3:0] _GEN_372; // @[StoreQueue.scala 75:25:@510.4]
  wire  _GEN_373; // @[StoreQueue.scala 75:25:@510.4]
  wire [3:0] _T_2002; // @[:@532.6]
  wire [3:0] _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_389; // @[StoreQueue.scala 76:20:@533.6]
  wire [3:0] _GEN_406; // @[StoreQueue.scala 75:25:@526.4]
  wire  _GEN_407; // @[StoreQueue.scala 75:25:@526.4]
  wire [3:0] _T_2020; // @[:@548.6]
  wire [3:0] _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_423; // @[StoreQueue.scala 76:20:@549.6]
  wire [3:0] _GEN_440; // @[StoreQueue.scala 75:25:@542.4]
  wire  _GEN_441; // @[StoreQueue.scala 75:25:@542.4]
  wire [3:0] _T_2038; // @[:@564.6]
  wire [3:0] _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_457; // @[StoreQueue.scala 76:20:@565.6]
  wire [3:0] _GEN_474; // @[StoreQueue.scala 75:25:@558.4]
  wire  _GEN_475; // @[StoreQueue.scala 75:25:@558.4]
  wire [3:0] _T_2056; // @[:@580.6]
  wire [3:0] _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_491; // @[StoreQueue.scala 76:20:@581.6]
  wire [3:0] _GEN_508; // @[StoreQueue.scala 75:25:@574.4]
  wire  _GEN_509; // @[StoreQueue.scala 75:25:@574.4]
  wire [3:0] _T_2074; // @[:@596.6]
  wire [3:0] _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_525; // @[StoreQueue.scala 76:20:@597.6]
  wire [3:0] _GEN_542; // @[StoreQueue.scala 75:25:@590.4]
  wire  _GEN_543; // @[StoreQueue.scala 75:25:@590.4]
  reg [3:0] previousLoadHead; // @[StoreQueue.scala 92:33:@606.4]
  reg [31:0] _RAND_146;
  wire [4:0] _T_2096; // @[util.scala 10:8:@615.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@616.6]
  wire [4:0] _T_2097; // @[util.scala 10:14:@616.6]
  wire [4:0] _GEN_1203; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2098; // @[StoreQueue.scala 96:56:@617.6]
  wire  _T_2099; // @[StoreQueue.scala 95:50:@618.6]
  wire  _T_2101; // @[StoreQueue.scala 95:35:@619.6]
  wire  _T_2103; // @[StoreQueue.scala 100:35:@627.8]
  wire  _T_2104; // @[StoreQueue.scala 100:87:@628.8]
  wire  _T_2105; // @[StoreQueue.scala 100:61:@629.8]
  wire  _T_2107; // @[StoreQueue.scala 102:35:@634.10]
  wire  _T_2108; // @[StoreQueue.scala 103:23:@635.10]
  wire  _T_2109; // @[StoreQueue.scala 103:75:@636.10]
  wire  _T_2110; // @[StoreQueue.scala 103:49:@637.10]
  wire  _T_2112; // @[StoreQueue.scala 103:9:@638.10]
  wire  _T_2113; // @[StoreQueue.scala 102:49:@639.10]
  wire  _GEN_560; // @[StoreQueue.scala 103:96:@640.10]
  wire  _GEN_561; // @[StoreQueue.scala 100:102:@630.8]
  wire  _GEN_562; // @[StoreQueue.scala 98:26:@623.6]
  wire  _GEN_563; // @[StoreQueue.scala 94:35:@608.4]
  wire [4:0] _T_2126; // @[util.scala 10:8:@651.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@652.6]
  wire [4:0] _T_2127; // @[util.scala 10:14:@652.6]
  wire  _T_2128; // @[StoreQueue.scala 96:56:@653.6]
  wire  _T_2129; // @[StoreQueue.scala 95:50:@654.6]
  wire  _T_2131; // @[StoreQueue.scala 95:35:@655.6]
  wire  _T_2133; // @[StoreQueue.scala 100:35:@663.8]
  wire  _T_2134; // @[StoreQueue.scala 100:87:@664.8]
  wire  _T_2135; // @[StoreQueue.scala 100:61:@665.8]
  wire  _T_2138; // @[StoreQueue.scala 103:23:@671.10]
  wire  _T_2139; // @[StoreQueue.scala 103:75:@672.10]
  wire  _T_2140; // @[StoreQueue.scala 103:49:@673.10]
  wire  _T_2142; // @[StoreQueue.scala 103:9:@674.10]
  wire  _T_2143; // @[StoreQueue.scala 102:49:@675.10]
  wire  _GEN_580; // @[StoreQueue.scala 103:96:@676.10]
  wire  _GEN_581; // @[StoreQueue.scala 100:102:@666.8]
  wire  _GEN_582; // @[StoreQueue.scala 98:26:@659.6]
  wire  _GEN_583; // @[StoreQueue.scala 94:35:@644.4]
  wire [4:0] _T_2156; // @[util.scala 10:8:@687.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@688.6]
  wire [4:0] _T_2157; // @[util.scala 10:14:@688.6]
  wire  _T_2158; // @[StoreQueue.scala 96:56:@689.6]
  wire  _T_2159; // @[StoreQueue.scala 95:50:@690.6]
  wire  _T_2161; // @[StoreQueue.scala 95:35:@691.6]
  wire  _T_2163; // @[StoreQueue.scala 100:35:@699.8]
  wire  _T_2164; // @[StoreQueue.scala 100:87:@700.8]
  wire  _T_2165; // @[StoreQueue.scala 100:61:@701.8]
  wire  _T_2168; // @[StoreQueue.scala 103:23:@707.10]
  wire  _T_2169; // @[StoreQueue.scala 103:75:@708.10]
  wire  _T_2170; // @[StoreQueue.scala 103:49:@709.10]
  wire  _T_2172; // @[StoreQueue.scala 103:9:@710.10]
  wire  _T_2173; // @[StoreQueue.scala 102:49:@711.10]
  wire  _GEN_600; // @[StoreQueue.scala 103:96:@712.10]
  wire  _GEN_601; // @[StoreQueue.scala 100:102:@702.8]
  wire  _GEN_602; // @[StoreQueue.scala 98:26:@695.6]
  wire  _GEN_603; // @[StoreQueue.scala 94:35:@680.4]
  wire [4:0] _T_2186; // @[util.scala 10:8:@723.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@724.6]
  wire [4:0] _T_2187; // @[util.scala 10:14:@724.6]
  wire  _T_2188; // @[StoreQueue.scala 96:56:@725.6]
  wire  _T_2189; // @[StoreQueue.scala 95:50:@726.6]
  wire  _T_2191; // @[StoreQueue.scala 95:35:@727.6]
  wire  _T_2193; // @[StoreQueue.scala 100:35:@735.8]
  wire  _T_2194; // @[StoreQueue.scala 100:87:@736.8]
  wire  _T_2195; // @[StoreQueue.scala 100:61:@737.8]
  wire  _T_2198; // @[StoreQueue.scala 103:23:@743.10]
  wire  _T_2199; // @[StoreQueue.scala 103:75:@744.10]
  wire  _T_2200; // @[StoreQueue.scala 103:49:@745.10]
  wire  _T_2202; // @[StoreQueue.scala 103:9:@746.10]
  wire  _T_2203; // @[StoreQueue.scala 102:49:@747.10]
  wire  _GEN_620; // @[StoreQueue.scala 103:96:@748.10]
  wire  _GEN_621; // @[StoreQueue.scala 100:102:@738.8]
  wire  _GEN_622; // @[StoreQueue.scala 98:26:@731.6]
  wire  _GEN_623; // @[StoreQueue.scala 94:35:@716.4]
  wire [4:0] _T_2216; // @[util.scala 10:8:@759.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@760.6]
  wire [4:0] _T_2217; // @[util.scala 10:14:@760.6]
  wire  _T_2218; // @[StoreQueue.scala 96:56:@761.6]
  wire  _T_2219; // @[StoreQueue.scala 95:50:@762.6]
  wire  _T_2221; // @[StoreQueue.scala 95:35:@763.6]
  wire  _T_2223; // @[StoreQueue.scala 100:35:@771.8]
  wire  _T_2224; // @[StoreQueue.scala 100:87:@772.8]
  wire  _T_2225; // @[StoreQueue.scala 100:61:@773.8]
  wire  _T_2228; // @[StoreQueue.scala 103:23:@779.10]
  wire  _T_2229; // @[StoreQueue.scala 103:75:@780.10]
  wire  _T_2230; // @[StoreQueue.scala 103:49:@781.10]
  wire  _T_2232; // @[StoreQueue.scala 103:9:@782.10]
  wire  _T_2233; // @[StoreQueue.scala 102:49:@783.10]
  wire  _GEN_640; // @[StoreQueue.scala 103:96:@784.10]
  wire  _GEN_641; // @[StoreQueue.scala 100:102:@774.8]
  wire  _GEN_642; // @[StoreQueue.scala 98:26:@767.6]
  wire  _GEN_643; // @[StoreQueue.scala 94:35:@752.4]
  wire [4:0] _T_2246; // @[util.scala 10:8:@795.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@796.6]
  wire [4:0] _T_2247; // @[util.scala 10:14:@796.6]
  wire  _T_2248; // @[StoreQueue.scala 96:56:@797.6]
  wire  _T_2249; // @[StoreQueue.scala 95:50:@798.6]
  wire  _T_2251; // @[StoreQueue.scala 95:35:@799.6]
  wire  _T_2253; // @[StoreQueue.scala 100:35:@807.8]
  wire  _T_2254; // @[StoreQueue.scala 100:87:@808.8]
  wire  _T_2255; // @[StoreQueue.scala 100:61:@809.8]
  wire  _T_2258; // @[StoreQueue.scala 103:23:@815.10]
  wire  _T_2259; // @[StoreQueue.scala 103:75:@816.10]
  wire  _T_2260; // @[StoreQueue.scala 103:49:@817.10]
  wire  _T_2262; // @[StoreQueue.scala 103:9:@818.10]
  wire  _T_2263; // @[StoreQueue.scala 102:49:@819.10]
  wire  _GEN_660; // @[StoreQueue.scala 103:96:@820.10]
  wire  _GEN_661; // @[StoreQueue.scala 100:102:@810.8]
  wire  _GEN_662; // @[StoreQueue.scala 98:26:@803.6]
  wire  _GEN_663; // @[StoreQueue.scala 94:35:@788.4]
  wire [4:0] _T_2276; // @[util.scala 10:8:@831.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@832.6]
  wire [4:0] _T_2277; // @[util.scala 10:14:@832.6]
  wire  _T_2278; // @[StoreQueue.scala 96:56:@833.6]
  wire  _T_2279; // @[StoreQueue.scala 95:50:@834.6]
  wire  _T_2281; // @[StoreQueue.scala 95:35:@835.6]
  wire  _T_2283; // @[StoreQueue.scala 100:35:@843.8]
  wire  _T_2284; // @[StoreQueue.scala 100:87:@844.8]
  wire  _T_2285; // @[StoreQueue.scala 100:61:@845.8]
  wire  _T_2288; // @[StoreQueue.scala 103:23:@851.10]
  wire  _T_2289; // @[StoreQueue.scala 103:75:@852.10]
  wire  _T_2290; // @[StoreQueue.scala 103:49:@853.10]
  wire  _T_2292; // @[StoreQueue.scala 103:9:@854.10]
  wire  _T_2293; // @[StoreQueue.scala 102:49:@855.10]
  wire  _GEN_680; // @[StoreQueue.scala 103:96:@856.10]
  wire  _GEN_681; // @[StoreQueue.scala 100:102:@846.8]
  wire  _GEN_682; // @[StoreQueue.scala 98:26:@839.6]
  wire  _GEN_683; // @[StoreQueue.scala 94:35:@824.4]
  wire [4:0] _T_2306; // @[util.scala 10:8:@867.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@868.6]
  wire [4:0] _T_2307; // @[util.scala 10:14:@868.6]
  wire  _T_2308; // @[StoreQueue.scala 96:56:@869.6]
  wire  _T_2309; // @[StoreQueue.scala 95:50:@870.6]
  wire  _T_2311; // @[StoreQueue.scala 95:35:@871.6]
  wire  _T_2313; // @[StoreQueue.scala 100:35:@879.8]
  wire  _T_2314; // @[StoreQueue.scala 100:87:@880.8]
  wire  _T_2315; // @[StoreQueue.scala 100:61:@881.8]
  wire  _T_2318; // @[StoreQueue.scala 103:23:@887.10]
  wire  _T_2319; // @[StoreQueue.scala 103:75:@888.10]
  wire  _T_2320; // @[StoreQueue.scala 103:49:@889.10]
  wire  _T_2322; // @[StoreQueue.scala 103:9:@890.10]
  wire  _T_2323; // @[StoreQueue.scala 102:49:@891.10]
  wire  _GEN_700; // @[StoreQueue.scala 103:96:@892.10]
  wire  _GEN_701; // @[StoreQueue.scala 100:102:@882.8]
  wire  _GEN_702; // @[StoreQueue.scala 98:26:@875.6]
  wire  _GEN_703; // @[StoreQueue.scala 94:35:@860.4]
  wire [4:0] _T_2336; // @[util.scala 10:8:@903.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@904.6]
  wire [4:0] _T_2337; // @[util.scala 10:14:@904.6]
  wire  _T_2338; // @[StoreQueue.scala 96:56:@905.6]
  wire  _T_2339; // @[StoreQueue.scala 95:50:@906.6]
  wire  _T_2341; // @[StoreQueue.scala 95:35:@907.6]
  wire  _T_2343; // @[StoreQueue.scala 100:35:@915.8]
  wire  _T_2344; // @[StoreQueue.scala 100:87:@916.8]
  wire  _T_2345; // @[StoreQueue.scala 100:61:@917.8]
  wire  _T_2348; // @[StoreQueue.scala 103:23:@923.10]
  wire  _T_2349; // @[StoreQueue.scala 103:75:@924.10]
  wire  _T_2350; // @[StoreQueue.scala 103:49:@925.10]
  wire  _T_2352; // @[StoreQueue.scala 103:9:@926.10]
  wire  _T_2353; // @[StoreQueue.scala 102:49:@927.10]
  wire  _GEN_720; // @[StoreQueue.scala 103:96:@928.10]
  wire  _GEN_721; // @[StoreQueue.scala 100:102:@918.8]
  wire  _GEN_722; // @[StoreQueue.scala 98:26:@911.6]
  wire  _GEN_723; // @[StoreQueue.scala 94:35:@896.4]
  wire [4:0] _T_2366; // @[util.scala 10:8:@939.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@940.6]
  wire [4:0] _T_2367; // @[util.scala 10:14:@940.6]
  wire  _T_2368; // @[StoreQueue.scala 96:56:@941.6]
  wire  _T_2369; // @[StoreQueue.scala 95:50:@942.6]
  wire  _T_2371; // @[StoreQueue.scala 95:35:@943.6]
  wire  _T_2373; // @[StoreQueue.scala 100:35:@951.8]
  wire  _T_2374; // @[StoreQueue.scala 100:87:@952.8]
  wire  _T_2375; // @[StoreQueue.scala 100:61:@953.8]
  wire  _T_2378; // @[StoreQueue.scala 103:23:@959.10]
  wire  _T_2379; // @[StoreQueue.scala 103:75:@960.10]
  wire  _T_2380; // @[StoreQueue.scala 103:49:@961.10]
  wire  _T_2382; // @[StoreQueue.scala 103:9:@962.10]
  wire  _T_2383; // @[StoreQueue.scala 102:49:@963.10]
  wire  _GEN_740; // @[StoreQueue.scala 103:96:@964.10]
  wire  _GEN_741; // @[StoreQueue.scala 100:102:@954.8]
  wire  _GEN_742; // @[StoreQueue.scala 98:26:@947.6]
  wire  _GEN_743; // @[StoreQueue.scala 94:35:@932.4]
  wire [4:0] _T_2396; // @[util.scala 10:8:@975.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@976.6]
  wire [4:0] _T_2397; // @[util.scala 10:14:@976.6]
  wire  _T_2398; // @[StoreQueue.scala 96:56:@977.6]
  wire  _T_2399; // @[StoreQueue.scala 95:50:@978.6]
  wire  _T_2401; // @[StoreQueue.scala 95:35:@979.6]
  wire  _T_2403; // @[StoreQueue.scala 100:35:@987.8]
  wire  _T_2404; // @[StoreQueue.scala 100:87:@988.8]
  wire  _T_2405; // @[StoreQueue.scala 100:61:@989.8]
  wire  _T_2408; // @[StoreQueue.scala 103:23:@995.10]
  wire  _T_2409; // @[StoreQueue.scala 103:75:@996.10]
  wire  _T_2410; // @[StoreQueue.scala 103:49:@997.10]
  wire  _T_2412; // @[StoreQueue.scala 103:9:@998.10]
  wire  _T_2413; // @[StoreQueue.scala 102:49:@999.10]
  wire  _GEN_760; // @[StoreQueue.scala 103:96:@1000.10]
  wire  _GEN_761; // @[StoreQueue.scala 100:102:@990.8]
  wire  _GEN_762; // @[StoreQueue.scala 98:26:@983.6]
  wire  _GEN_763; // @[StoreQueue.scala 94:35:@968.4]
  wire [4:0] _T_2426; // @[util.scala 10:8:@1011.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@1012.6]
  wire [4:0] _T_2427; // @[util.scala 10:14:@1012.6]
  wire  _T_2428; // @[StoreQueue.scala 96:56:@1013.6]
  wire  _T_2429; // @[StoreQueue.scala 95:50:@1014.6]
  wire  _T_2431; // @[StoreQueue.scala 95:35:@1015.6]
  wire  _T_2433; // @[StoreQueue.scala 100:35:@1023.8]
  wire  _T_2434; // @[StoreQueue.scala 100:87:@1024.8]
  wire  _T_2435; // @[StoreQueue.scala 100:61:@1025.8]
  wire  _T_2438; // @[StoreQueue.scala 103:23:@1031.10]
  wire  _T_2439; // @[StoreQueue.scala 103:75:@1032.10]
  wire  _T_2440; // @[StoreQueue.scala 103:49:@1033.10]
  wire  _T_2442; // @[StoreQueue.scala 103:9:@1034.10]
  wire  _T_2443; // @[StoreQueue.scala 102:49:@1035.10]
  wire  _GEN_780; // @[StoreQueue.scala 103:96:@1036.10]
  wire  _GEN_781; // @[StoreQueue.scala 100:102:@1026.8]
  wire  _GEN_782; // @[StoreQueue.scala 98:26:@1019.6]
  wire  _GEN_783; // @[StoreQueue.scala 94:35:@1004.4]
  wire [4:0] _T_2456; // @[util.scala 10:8:@1047.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@1048.6]
  wire [4:0] _T_2457; // @[util.scala 10:14:@1048.6]
  wire  _T_2458; // @[StoreQueue.scala 96:56:@1049.6]
  wire  _T_2459; // @[StoreQueue.scala 95:50:@1050.6]
  wire  _T_2461; // @[StoreQueue.scala 95:35:@1051.6]
  wire  _T_2463; // @[StoreQueue.scala 100:35:@1059.8]
  wire  _T_2464; // @[StoreQueue.scala 100:87:@1060.8]
  wire  _T_2465; // @[StoreQueue.scala 100:61:@1061.8]
  wire  _T_2468; // @[StoreQueue.scala 103:23:@1067.10]
  wire  _T_2469; // @[StoreQueue.scala 103:75:@1068.10]
  wire  _T_2470; // @[StoreQueue.scala 103:49:@1069.10]
  wire  _T_2472; // @[StoreQueue.scala 103:9:@1070.10]
  wire  _T_2473; // @[StoreQueue.scala 102:49:@1071.10]
  wire  _GEN_800; // @[StoreQueue.scala 103:96:@1072.10]
  wire  _GEN_801; // @[StoreQueue.scala 100:102:@1062.8]
  wire  _GEN_802; // @[StoreQueue.scala 98:26:@1055.6]
  wire  _GEN_803; // @[StoreQueue.scala 94:35:@1040.4]
  wire [4:0] _T_2486; // @[util.scala 10:8:@1083.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@1084.6]
  wire [4:0] _T_2487; // @[util.scala 10:14:@1084.6]
  wire  _T_2488; // @[StoreQueue.scala 96:56:@1085.6]
  wire  _T_2489; // @[StoreQueue.scala 95:50:@1086.6]
  wire  _T_2491; // @[StoreQueue.scala 95:35:@1087.6]
  wire  _T_2493; // @[StoreQueue.scala 100:35:@1095.8]
  wire  _T_2494; // @[StoreQueue.scala 100:87:@1096.8]
  wire  _T_2495; // @[StoreQueue.scala 100:61:@1097.8]
  wire  _T_2498; // @[StoreQueue.scala 103:23:@1103.10]
  wire  _T_2499; // @[StoreQueue.scala 103:75:@1104.10]
  wire  _T_2500; // @[StoreQueue.scala 103:49:@1105.10]
  wire  _T_2502; // @[StoreQueue.scala 103:9:@1106.10]
  wire  _T_2503; // @[StoreQueue.scala 102:49:@1107.10]
  wire  _GEN_820; // @[StoreQueue.scala 103:96:@1108.10]
  wire  _GEN_821; // @[StoreQueue.scala 100:102:@1098.8]
  wire  _GEN_822; // @[StoreQueue.scala 98:26:@1091.6]
  wire  _GEN_823; // @[StoreQueue.scala 94:35:@1076.4]
  wire [4:0] _T_2516; // @[util.scala 10:8:@1119.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@1120.6]
  wire [4:0] _T_2517; // @[util.scala 10:14:@1120.6]
  wire  _T_2518; // @[StoreQueue.scala 96:56:@1121.6]
  wire  _T_2519; // @[StoreQueue.scala 95:50:@1122.6]
  wire  _T_2521; // @[StoreQueue.scala 95:35:@1123.6]
  wire  _T_2523; // @[StoreQueue.scala 100:35:@1131.8]
  wire  _T_2524; // @[StoreQueue.scala 100:87:@1132.8]
  wire  _T_2525; // @[StoreQueue.scala 100:61:@1133.8]
  wire  _T_2528; // @[StoreQueue.scala 103:23:@1139.10]
  wire  _T_2529; // @[StoreQueue.scala 103:75:@1140.10]
  wire  _T_2530; // @[StoreQueue.scala 103:49:@1141.10]
  wire  _T_2532; // @[StoreQueue.scala 103:9:@1142.10]
  wire  _T_2533; // @[StoreQueue.scala 102:49:@1143.10]
  wire  _GEN_840; // @[StoreQueue.scala 103:96:@1144.10]
  wire  _GEN_841; // @[StoreQueue.scala 100:102:@1134.8]
  wire  _GEN_842; // @[StoreQueue.scala 98:26:@1127.6]
  wire  _GEN_843; // @[StoreQueue.scala 94:35:@1112.4]
  wire [4:0] _T_2546; // @[util.scala 10:8:@1155.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@1156.6]
  wire [4:0] _T_2547; // @[util.scala 10:14:@1156.6]
  wire  _T_2548; // @[StoreQueue.scala 96:56:@1157.6]
  wire  _T_2549; // @[StoreQueue.scala 95:50:@1158.6]
  wire  _T_2551; // @[StoreQueue.scala 95:35:@1159.6]
  wire  _T_2553; // @[StoreQueue.scala 100:35:@1167.8]
  wire  _T_2554; // @[StoreQueue.scala 100:87:@1168.8]
  wire  _T_2555; // @[StoreQueue.scala 100:61:@1169.8]
  wire  _T_2558; // @[StoreQueue.scala 103:23:@1175.10]
  wire  _T_2559; // @[StoreQueue.scala 103:75:@1176.10]
  wire  _T_2560; // @[StoreQueue.scala 103:49:@1177.10]
  wire  _T_2562; // @[StoreQueue.scala 103:9:@1178.10]
  wire  _T_2563; // @[StoreQueue.scala 102:49:@1179.10]
  wire  _GEN_860; // @[StoreQueue.scala 103:96:@1180.10]
  wire  _GEN_861; // @[StoreQueue.scala 100:102:@1170.8]
  wire  _GEN_862; // @[StoreQueue.scala 98:26:@1163.6]
  wire  _GEN_863; // @[StoreQueue.scala 94:35:@1148.4]
  wire  _T_2565; // @[StoreQueue.scala 119:103:@1184.4]
  wire  _T_2567; // @[StoreQueue.scala 120:17:@1185.4]
  wire  _T_2569; // @[StoreQueue.scala 120:35:@1186.4]
  wire  _T_2570; // @[StoreQueue.scala 120:26:@1187.4]
  wire  _T_2572; // @[StoreQueue.scala 120:50:@1188.4]
  wire  _T_2574; // @[StoreQueue.scala 120:81:@1189.4]
  wire  _T_2576; // @[StoreQueue.scala 120:99:@1190.4]
  wire  _T_2577; // @[StoreQueue.scala 120:90:@1191.4]
  wire  _T_2579; // @[StoreQueue.scala 120:67:@1192.4]
  wire  _T_2580; // @[StoreQueue.scala 120:64:@1193.4]
  wire  validEntriesInLoadQ_0; // @[StoreQueue.scala 119:90:@1194.4]
  wire  _T_2584; // @[StoreQueue.scala 120:17:@1196.4]
  wire  _T_2586; // @[StoreQueue.scala 120:35:@1197.4]
  wire  _T_2587; // @[StoreQueue.scala 120:26:@1198.4]
  wire  _T_2591; // @[StoreQueue.scala 120:81:@1200.4]
  wire  _T_2593; // @[StoreQueue.scala 120:99:@1201.4]
  wire  _T_2594; // @[StoreQueue.scala 120:90:@1202.4]
  wire  _T_2596; // @[StoreQueue.scala 120:67:@1203.4]
  wire  _T_2597; // @[StoreQueue.scala 120:64:@1204.4]
  wire  validEntriesInLoadQ_1; // @[StoreQueue.scala 119:90:@1205.4]
  wire  _T_2601; // @[StoreQueue.scala 120:17:@1207.4]
  wire  _T_2603; // @[StoreQueue.scala 120:35:@1208.4]
  wire  _T_2604; // @[StoreQueue.scala 120:26:@1209.4]
  wire  _T_2608; // @[StoreQueue.scala 120:81:@1211.4]
  wire  _T_2610; // @[StoreQueue.scala 120:99:@1212.4]
  wire  _T_2611; // @[StoreQueue.scala 120:90:@1213.4]
  wire  _T_2613; // @[StoreQueue.scala 120:67:@1214.4]
  wire  _T_2614; // @[StoreQueue.scala 120:64:@1215.4]
  wire  validEntriesInLoadQ_2; // @[StoreQueue.scala 119:90:@1216.4]
  wire  _T_2618; // @[StoreQueue.scala 120:17:@1218.4]
  wire  _T_2620; // @[StoreQueue.scala 120:35:@1219.4]
  wire  _T_2621; // @[StoreQueue.scala 120:26:@1220.4]
  wire  _T_2625; // @[StoreQueue.scala 120:81:@1222.4]
  wire  _T_2627; // @[StoreQueue.scala 120:99:@1223.4]
  wire  _T_2628; // @[StoreQueue.scala 120:90:@1224.4]
  wire  _T_2630; // @[StoreQueue.scala 120:67:@1225.4]
  wire  _T_2631; // @[StoreQueue.scala 120:64:@1226.4]
  wire  validEntriesInLoadQ_3; // @[StoreQueue.scala 119:90:@1227.4]
  wire  _T_2635; // @[StoreQueue.scala 120:17:@1229.4]
  wire  _T_2637; // @[StoreQueue.scala 120:35:@1230.4]
  wire  _T_2638; // @[StoreQueue.scala 120:26:@1231.4]
  wire  _T_2642; // @[StoreQueue.scala 120:81:@1233.4]
  wire  _T_2644; // @[StoreQueue.scala 120:99:@1234.4]
  wire  _T_2645; // @[StoreQueue.scala 120:90:@1235.4]
  wire  _T_2647; // @[StoreQueue.scala 120:67:@1236.4]
  wire  _T_2648; // @[StoreQueue.scala 120:64:@1237.4]
  wire  validEntriesInLoadQ_4; // @[StoreQueue.scala 119:90:@1238.4]
  wire  _T_2652; // @[StoreQueue.scala 120:17:@1240.4]
  wire  _T_2654; // @[StoreQueue.scala 120:35:@1241.4]
  wire  _T_2655; // @[StoreQueue.scala 120:26:@1242.4]
  wire  _T_2659; // @[StoreQueue.scala 120:81:@1244.4]
  wire  _T_2661; // @[StoreQueue.scala 120:99:@1245.4]
  wire  _T_2662; // @[StoreQueue.scala 120:90:@1246.4]
  wire  _T_2664; // @[StoreQueue.scala 120:67:@1247.4]
  wire  _T_2665; // @[StoreQueue.scala 120:64:@1248.4]
  wire  validEntriesInLoadQ_5; // @[StoreQueue.scala 119:90:@1249.4]
  wire  _T_2669; // @[StoreQueue.scala 120:17:@1251.4]
  wire  _T_2671; // @[StoreQueue.scala 120:35:@1252.4]
  wire  _T_2672; // @[StoreQueue.scala 120:26:@1253.4]
  wire  _T_2676; // @[StoreQueue.scala 120:81:@1255.4]
  wire  _T_2678; // @[StoreQueue.scala 120:99:@1256.4]
  wire  _T_2679; // @[StoreQueue.scala 120:90:@1257.4]
  wire  _T_2681; // @[StoreQueue.scala 120:67:@1258.4]
  wire  _T_2682; // @[StoreQueue.scala 120:64:@1259.4]
  wire  validEntriesInLoadQ_6; // @[StoreQueue.scala 119:90:@1260.4]
  wire  _T_2686; // @[StoreQueue.scala 120:17:@1262.4]
  wire  _T_2688; // @[StoreQueue.scala 120:35:@1263.4]
  wire  _T_2689; // @[StoreQueue.scala 120:26:@1264.4]
  wire  _T_2693; // @[StoreQueue.scala 120:81:@1266.4]
  wire  _T_2695; // @[StoreQueue.scala 120:99:@1267.4]
  wire  _T_2696; // @[StoreQueue.scala 120:90:@1268.4]
  wire  _T_2698; // @[StoreQueue.scala 120:67:@1269.4]
  wire  _T_2699; // @[StoreQueue.scala 120:64:@1270.4]
  wire  validEntriesInLoadQ_7; // @[StoreQueue.scala 119:90:@1271.4]
  wire  _T_2703; // @[StoreQueue.scala 120:17:@1273.4]
  wire  _T_2705; // @[StoreQueue.scala 120:35:@1274.4]
  wire  _T_2706; // @[StoreQueue.scala 120:26:@1275.4]
  wire  _T_2710; // @[StoreQueue.scala 120:81:@1277.4]
  wire  _T_2712; // @[StoreQueue.scala 120:99:@1278.4]
  wire  _T_2713; // @[StoreQueue.scala 120:90:@1279.4]
  wire  _T_2715; // @[StoreQueue.scala 120:67:@1280.4]
  wire  _T_2716; // @[StoreQueue.scala 120:64:@1281.4]
  wire  validEntriesInLoadQ_8; // @[StoreQueue.scala 119:90:@1282.4]
  wire  _T_2720; // @[StoreQueue.scala 120:17:@1284.4]
  wire  _T_2722; // @[StoreQueue.scala 120:35:@1285.4]
  wire  _T_2723; // @[StoreQueue.scala 120:26:@1286.4]
  wire  _T_2727; // @[StoreQueue.scala 120:81:@1288.4]
  wire  _T_2729; // @[StoreQueue.scala 120:99:@1289.4]
  wire  _T_2730; // @[StoreQueue.scala 120:90:@1290.4]
  wire  _T_2732; // @[StoreQueue.scala 120:67:@1291.4]
  wire  _T_2733; // @[StoreQueue.scala 120:64:@1292.4]
  wire  validEntriesInLoadQ_9; // @[StoreQueue.scala 119:90:@1293.4]
  wire  _T_2737; // @[StoreQueue.scala 120:17:@1295.4]
  wire  _T_2739; // @[StoreQueue.scala 120:35:@1296.4]
  wire  _T_2740; // @[StoreQueue.scala 120:26:@1297.4]
  wire  _T_2744; // @[StoreQueue.scala 120:81:@1299.4]
  wire  _T_2746; // @[StoreQueue.scala 120:99:@1300.4]
  wire  _T_2747; // @[StoreQueue.scala 120:90:@1301.4]
  wire  _T_2749; // @[StoreQueue.scala 120:67:@1302.4]
  wire  _T_2750; // @[StoreQueue.scala 120:64:@1303.4]
  wire  validEntriesInLoadQ_10; // @[StoreQueue.scala 119:90:@1304.4]
  wire  _T_2754; // @[StoreQueue.scala 120:17:@1306.4]
  wire  _T_2756; // @[StoreQueue.scala 120:35:@1307.4]
  wire  _T_2757; // @[StoreQueue.scala 120:26:@1308.4]
  wire  _T_2761; // @[StoreQueue.scala 120:81:@1310.4]
  wire  _T_2763; // @[StoreQueue.scala 120:99:@1311.4]
  wire  _T_2764; // @[StoreQueue.scala 120:90:@1312.4]
  wire  _T_2766; // @[StoreQueue.scala 120:67:@1313.4]
  wire  _T_2767; // @[StoreQueue.scala 120:64:@1314.4]
  wire  validEntriesInLoadQ_11; // @[StoreQueue.scala 119:90:@1315.4]
  wire  _T_2771; // @[StoreQueue.scala 120:17:@1317.4]
  wire  _T_2773; // @[StoreQueue.scala 120:35:@1318.4]
  wire  _T_2774; // @[StoreQueue.scala 120:26:@1319.4]
  wire  _T_2778; // @[StoreQueue.scala 120:81:@1321.4]
  wire  _T_2780; // @[StoreQueue.scala 120:99:@1322.4]
  wire  _T_2781; // @[StoreQueue.scala 120:90:@1323.4]
  wire  _T_2783; // @[StoreQueue.scala 120:67:@1324.4]
  wire  _T_2784; // @[StoreQueue.scala 120:64:@1325.4]
  wire  validEntriesInLoadQ_12; // @[StoreQueue.scala 119:90:@1326.4]
  wire  _T_2788; // @[StoreQueue.scala 120:17:@1328.4]
  wire  _T_2790; // @[StoreQueue.scala 120:35:@1329.4]
  wire  _T_2791; // @[StoreQueue.scala 120:26:@1330.4]
  wire  _T_2795; // @[StoreQueue.scala 120:81:@1332.4]
  wire  _T_2797; // @[StoreQueue.scala 120:99:@1333.4]
  wire  _T_2798; // @[StoreQueue.scala 120:90:@1334.4]
  wire  _T_2800; // @[StoreQueue.scala 120:67:@1335.4]
  wire  _T_2801; // @[StoreQueue.scala 120:64:@1336.4]
  wire  validEntriesInLoadQ_13; // @[StoreQueue.scala 119:90:@1337.4]
  wire  _T_2805; // @[StoreQueue.scala 120:17:@1339.4]
  wire  _T_2807; // @[StoreQueue.scala 120:35:@1340.4]
  wire  _T_2808; // @[StoreQueue.scala 120:26:@1341.4]
  wire  _T_2812; // @[StoreQueue.scala 120:81:@1343.4]
  wire  _T_2814; // @[StoreQueue.scala 120:99:@1344.4]
  wire  _T_2815; // @[StoreQueue.scala 120:90:@1345.4]
  wire  _T_2817; // @[StoreQueue.scala 120:67:@1346.4]
  wire  _T_2818; // @[StoreQueue.scala 120:64:@1347.4]
  wire  validEntriesInLoadQ_14; // @[StoreQueue.scala 119:90:@1348.4]
  wire  validEntriesInLoadQ_15; // @[StoreQueue.scala 119:90:@1359.4]
  wire [3:0] _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  wire [3:0] _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  wire  _T_2861; // @[StoreQueue.scala 126:96:@1377.4]
  wire  loadsToCheck_0; // @[StoreQueue.scala 126:83:@1385.4]
  wire  _T_2891; // @[StoreQueue.scala 127:37:@1388.4]
  wire  _T_2892; // @[StoreQueue.scala 127:28:@1389.4]
  wire  _T_2897; // @[StoreQueue.scala 127:71:@1390.4]
  wire  _T_2900; // @[StoreQueue.scala 127:79:@1392.4]
  wire  _T_2902; // @[StoreQueue.scala 127:55:@1393.4]
  wire  loadsToCheck_1; // @[StoreQueue.scala 126:83:@1394.4]
  wire  _T_2914; // @[StoreQueue.scala 127:37:@1397.4]
  wire  _T_2915; // @[StoreQueue.scala 127:28:@1398.4]
  wire  _T_2920; // @[StoreQueue.scala 127:71:@1399.4]
  wire  _T_2923; // @[StoreQueue.scala 127:79:@1401.4]
  wire  _T_2925; // @[StoreQueue.scala 127:55:@1402.4]
  wire  loadsToCheck_2; // @[StoreQueue.scala 126:83:@1403.4]
  wire  _T_2937; // @[StoreQueue.scala 127:37:@1406.4]
  wire  _T_2938; // @[StoreQueue.scala 127:28:@1407.4]
  wire  _T_2943; // @[StoreQueue.scala 127:71:@1408.4]
  wire  _T_2946; // @[StoreQueue.scala 127:79:@1410.4]
  wire  _T_2948; // @[StoreQueue.scala 127:55:@1411.4]
  wire  loadsToCheck_3; // @[StoreQueue.scala 126:83:@1412.4]
  wire  _T_2960; // @[StoreQueue.scala 127:37:@1415.4]
  wire  _T_2961; // @[StoreQueue.scala 127:28:@1416.4]
  wire  _T_2966; // @[StoreQueue.scala 127:71:@1417.4]
  wire  _T_2969; // @[StoreQueue.scala 127:79:@1419.4]
  wire  _T_2971; // @[StoreQueue.scala 127:55:@1420.4]
  wire  loadsToCheck_4; // @[StoreQueue.scala 126:83:@1421.4]
  wire  _T_2983; // @[StoreQueue.scala 127:37:@1424.4]
  wire  _T_2984; // @[StoreQueue.scala 127:28:@1425.4]
  wire  _T_2989; // @[StoreQueue.scala 127:71:@1426.4]
  wire  _T_2992; // @[StoreQueue.scala 127:79:@1428.4]
  wire  _T_2994; // @[StoreQueue.scala 127:55:@1429.4]
  wire  loadsToCheck_5; // @[StoreQueue.scala 126:83:@1430.4]
  wire  _T_3006; // @[StoreQueue.scala 127:37:@1433.4]
  wire  _T_3007; // @[StoreQueue.scala 127:28:@1434.4]
  wire  _T_3012; // @[StoreQueue.scala 127:71:@1435.4]
  wire  _T_3015; // @[StoreQueue.scala 127:79:@1437.4]
  wire  _T_3017; // @[StoreQueue.scala 127:55:@1438.4]
  wire  loadsToCheck_6; // @[StoreQueue.scala 126:83:@1439.4]
  wire  _T_3029; // @[StoreQueue.scala 127:37:@1442.4]
  wire  _T_3030; // @[StoreQueue.scala 127:28:@1443.4]
  wire  _T_3035; // @[StoreQueue.scala 127:71:@1444.4]
  wire  _T_3038; // @[StoreQueue.scala 127:79:@1446.4]
  wire  _T_3040; // @[StoreQueue.scala 127:55:@1447.4]
  wire  loadsToCheck_7; // @[StoreQueue.scala 126:83:@1448.4]
  wire  _T_3052; // @[StoreQueue.scala 127:37:@1451.4]
  wire  _T_3053; // @[StoreQueue.scala 127:28:@1452.4]
  wire  _T_3058; // @[StoreQueue.scala 127:71:@1453.4]
  wire  _T_3061; // @[StoreQueue.scala 127:79:@1455.4]
  wire  _T_3063; // @[StoreQueue.scala 127:55:@1456.4]
  wire  loadsToCheck_8; // @[StoreQueue.scala 126:83:@1457.4]
  wire  _T_3075; // @[StoreQueue.scala 127:37:@1460.4]
  wire  _T_3076; // @[StoreQueue.scala 127:28:@1461.4]
  wire  _T_3081; // @[StoreQueue.scala 127:71:@1462.4]
  wire  _T_3084; // @[StoreQueue.scala 127:79:@1464.4]
  wire  _T_3086; // @[StoreQueue.scala 127:55:@1465.4]
  wire  loadsToCheck_9; // @[StoreQueue.scala 126:83:@1466.4]
  wire  _T_3098; // @[StoreQueue.scala 127:37:@1469.4]
  wire  _T_3099; // @[StoreQueue.scala 127:28:@1470.4]
  wire  _T_3104; // @[StoreQueue.scala 127:71:@1471.4]
  wire  _T_3107; // @[StoreQueue.scala 127:79:@1473.4]
  wire  _T_3109; // @[StoreQueue.scala 127:55:@1474.4]
  wire  loadsToCheck_10; // @[StoreQueue.scala 126:83:@1475.4]
  wire  _T_3121; // @[StoreQueue.scala 127:37:@1478.4]
  wire  _T_3122; // @[StoreQueue.scala 127:28:@1479.4]
  wire  _T_3127; // @[StoreQueue.scala 127:71:@1480.4]
  wire  _T_3130; // @[StoreQueue.scala 127:79:@1482.4]
  wire  _T_3132; // @[StoreQueue.scala 127:55:@1483.4]
  wire  loadsToCheck_11; // @[StoreQueue.scala 126:83:@1484.4]
  wire  _T_3144; // @[StoreQueue.scala 127:37:@1487.4]
  wire  _T_3145; // @[StoreQueue.scala 127:28:@1488.4]
  wire  _T_3150; // @[StoreQueue.scala 127:71:@1489.4]
  wire  _T_3153; // @[StoreQueue.scala 127:79:@1491.4]
  wire  _T_3155; // @[StoreQueue.scala 127:55:@1492.4]
  wire  loadsToCheck_12; // @[StoreQueue.scala 126:83:@1493.4]
  wire  _T_3167; // @[StoreQueue.scala 127:37:@1496.4]
  wire  _T_3168; // @[StoreQueue.scala 127:28:@1497.4]
  wire  _T_3173; // @[StoreQueue.scala 127:71:@1498.4]
  wire  _T_3176; // @[StoreQueue.scala 127:79:@1500.4]
  wire  _T_3178; // @[StoreQueue.scala 127:55:@1501.4]
  wire  loadsToCheck_13; // @[StoreQueue.scala 126:83:@1502.4]
  wire  _T_3190; // @[StoreQueue.scala 127:37:@1505.4]
  wire  _T_3191; // @[StoreQueue.scala 127:28:@1506.4]
  wire  _T_3196; // @[StoreQueue.scala 127:71:@1507.4]
  wire  _T_3199; // @[StoreQueue.scala 127:79:@1509.4]
  wire  _T_3201; // @[StoreQueue.scala 127:55:@1510.4]
  wire  loadsToCheck_14; // @[StoreQueue.scala 126:83:@1511.4]
  wire  _T_3213; // @[StoreQueue.scala 127:37:@1514.4]
  wire  loadsToCheck_15; // @[StoreQueue.scala 126:83:@1520.4]
  wire  _T_3247; // @[StoreQueue.scala 133:16:@1538.4]
  wire  _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  wire  entriesToCheck_0; // @[StoreQueue.scala 133:24:@1539.4]
  wire  _T_3252; // @[StoreQueue.scala 133:16:@1540.4]
  wire  entriesToCheck_1; // @[StoreQueue.scala 133:24:@1541.4]
  wire  _T_3257; // @[StoreQueue.scala 133:16:@1542.4]
  wire  entriesToCheck_2; // @[StoreQueue.scala 133:24:@1543.4]
  wire  _T_3262; // @[StoreQueue.scala 133:16:@1544.4]
  wire  entriesToCheck_3; // @[StoreQueue.scala 133:24:@1545.4]
  wire  _T_3267; // @[StoreQueue.scala 133:16:@1546.4]
  wire  entriesToCheck_4; // @[StoreQueue.scala 133:24:@1547.4]
  wire  _T_3272; // @[StoreQueue.scala 133:16:@1548.4]
  wire  entriesToCheck_5; // @[StoreQueue.scala 133:24:@1549.4]
  wire  _T_3277; // @[StoreQueue.scala 133:16:@1550.4]
  wire  entriesToCheck_6; // @[StoreQueue.scala 133:24:@1551.4]
  wire  _T_3282; // @[StoreQueue.scala 133:16:@1552.4]
  wire  entriesToCheck_7; // @[StoreQueue.scala 133:24:@1553.4]
  wire  _T_3287; // @[StoreQueue.scala 133:16:@1554.4]
  wire  entriesToCheck_8; // @[StoreQueue.scala 133:24:@1555.4]
  wire  _T_3292; // @[StoreQueue.scala 133:16:@1556.4]
  wire  entriesToCheck_9; // @[StoreQueue.scala 133:24:@1557.4]
  wire  _T_3297; // @[StoreQueue.scala 133:16:@1558.4]
  wire  entriesToCheck_10; // @[StoreQueue.scala 133:24:@1559.4]
  wire  _T_3302; // @[StoreQueue.scala 133:16:@1560.4]
  wire  entriesToCheck_11; // @[StoreQueue.scala 133:24:@1561.4]
  wire  _T_3307; // @[StoreQueue.scala 133:16:@1562.4]
  wire  entriesToCheck_12; // @[StoreQueue.scala 133:24:@1563.4]
  wire  _T_3312; // @[StoreQueue.scala 133:16:@1564.4]
  wire  entriesToCheck_13; // @[StoreQueue.scala 133:24:@1565.4]
  wire  _T_3317; // @[StoreQueue.scala 133:16:@1566.4]
  wire  entriesToCheck_14; // @[StoreQueue.scala 133:24:@1567.4]
  wire  _T_3322; // @[StoreQueue.scala 133:16:@1568.4]
  wire  entriesToCheck_15; // @[StoreQueue.scala 133:24:@1569.4]
  wire  _T_3370; // @[StoreQueue.scala 140:34:@1588.4]
  wire  _T_3371; // @[StoreQueue.scala 140:64:@1589.4]
  wire [31:0] _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  wire [31:0] _GEN_911; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3375; // @[StoreQueue.scala 141:51:@1590.4]
  wire  _T_3376; // @[StoreQueue.scala 141:36:@1591.4]
  wire  noConflicts_0; // @[StoreQueue.scala 140:95:@1592.4]
  wire  _T_3379; // @[StoreQueue.scala 140:34:@1594.4]
  wire  _T_3380; // @[StoreQueue.scala 140:64:@1595.4]
  wire  _T_3384; // @[StoreQueue.scala 141:51:@1596.4]
  wire  _T_3385; // @[StoreQueue.scala 141:36:@1597.4]
  wire  noConflicts_1; // @[StoreQueue.scala 140:95:@1598.4]
  wire  _T_3388; // @[StoreQueue.scala 140:34:@1600.4]
  wire  _T_3389; // @[StoreQueue.scala 140:64:@1601.4]
  wire  _T_3393; // @[StoreQueue.scala 141:51:@1602.4]
  wire  _T_3394; // @[StoreQueue.scala 141:36:@1603.4]
  wire  noConflicts_2; // @[StoreQueue.scala 140:95:@1604.4]
  wire  _T_3397; // @[StoreQueue.scala 140:34:@1606.4]
  wire  _T_3398; // @[StoreQueue.scala 140:64:@1607.4]
  wire  _T_3402; // @[StoreQueue.scala 141:51:@1608.4]
  wire  _T_3403; // @[StoreQueue.scala 141:36:@1609.4]
  wire  noConflicts_3; // @[StoreQueue.scala 140:95:@1610.4]
  wire  _T_3406; // @[StoreQueue.scala 140:34:@1612.4]
  wire  _T_3407; // @[StoreQueue.scala 140:64:@1613.4]
  wire  _T_3411; // @[StoreQueue.scala 141:51:@1614.4]
  wire  _T_3412; // @[StoreQueue.scala 141:36:@1615.4]
  wire  noConflicts_4; // @[StoreQueue.scala 140:95:@1616.4]
  wire  _T_3415; // @[StoreQueue.scala 140:34:@1618.4]
  wire  _T_3416; // @[StoreQueue.scala 140:64:@1619.4]
  wire  _T_3420; // @[StoreQueue.scala 141:51:@1620.4]
  wire  _T_3421; // @[StoreQueue.scala 141:36:@1621.4]
  wire  noConflicts_5; // @[StoreQueue.scala 140:95:@1622.4]
  wire  _T_3424; // @[StoreQueue.scala 140:34:@1624.4]
  wire  _T_3425; // @[StoreQueue.scala 140:64:@1625.4]
  wire  _T_3429; // @[StoreQueue.scala 141:51:@1626.4]
  wire  _T_3430; // @[StoreQueue.scala 141:36:@1627.4]
  wire  noConflicts_6; // @[StoreQueue.scala 140:95:@1628.4]
  wire  _T_3433; // @[StoreQueue.scala 140:34:@1630.4]
  wire  _T_3434; // @[StoreQueue.scala 140:64:@1631.4]
  wire  _T_3438; // @[StoreQueue.scala 141:51:@1632.4]
  wire  _T_3439; // @[StoreQueue.scala 141:36:@1633.4]
  wire  noConflicts_7; // @[StoreQueue.scala 140:95:@1634.4]
  wire  _T_3442; // @[StoreQueue.scala 140:34:@1636.4]
  wire  _T_3443; // @[StoreQueue.scala 140:64:@1637.4]
  wire  _T_3447; // @[StoreQueue.scala 141:51:@1638.4]
  wire  _T_3448; // @[StoreQueue.scala 141:36:@1639.4]
  wire  noConflicts_8; // @[StoreQueue.scala 140:95:@1640.4]
  wire  _T_3451; // @[StoreQueue.scala 140:34:@1642.4]
  wire  _T_3452; // @[StoreQueue.scala 140:64:@1643.4]
  wire  _T_3456; // @[StoreQueue.scala 141:51:@1644.4]
  wire  _T_3457; // @[StoreQueue.scala 141:36:@1645.4]
  wire  noConflicts_9; // @[StoreQueue.scala 140:95:@1646.4]
  wire  _T_3460; // @[StoreQueue.scala 140:34:@1648.4]
  wire  _T_3461; // @[StoreQueue.scala 140:64:@1649.4]
  wire  _T_3465; // @[StoreQueue.scala 141:51:@1650.4]
  wire  _T_3466; // @[StoreQueue.scala 141:36:@1651.4]
  wire  noConflicts_10; // @[StoreQueue.scala 140:95:@1652.4]
  wire  _T_3469; // @[StoreQueue.scala 140:34:@1654.4]
  wire  _T_3470; // @[StoreQueue.scala 140:64:@1655.4]
  wire  _T_3474; // @[StoreQueue.scala 141:51:@1656.4]
  wire  _T_3475; // @[StoreQueue.scala 141:36:@1657.4]
  wire  noConflicts_11; // @[StoreQueue.scala 140:95:@1658.4]
  wire  _T_3478; // @[StoreQueue.scala 140:34:@1660.4]
  wire  _T_3479; // @[StoreQueue.scala 140:64:@1661.4]
  wire  _T_3483; // @[StoreQueue.scala 141:51:@1662.4]
  wire  _T_3484; // @[StoreQueue.scala 141:36:@1663.4]
  wire  noConflicts_12; // @[StoreQueue.scala 140:95:@1664.4]
  wire  _T_3487; // @[StoreQueue.scala 140:34:@1666.4]
  wire  _T_3488; // @[StoreQueue.scala 140:64:@1667.4]
  wire  _T_3492; // @[StoreQueue.scala 141:51:@1668.4]
  wire  _T_3493; // @[StoreQueue.scala 141:36:@1669.4]
  wire  noConflicts_13; // @[StoreQueue.scala 140:95:@1670.4]
  wire  _T_3496; // @[StoreQueue.scala 140:34:@1672.4]
  wire  _T_3497; // @[StoreQueue.scala 140:64:@1673.4]
  wire  _T_3501; // @[StoreQueue.scala 141:51:@1674.4]
  wire  _T_3502; // @[StoreQueue.scala 141:36:@1675.4]
  wire  noConflicts_14; // @[StoreQueue.scala 140:95:@1676.4]
  wire  _T_3505; // @[StoreQueue.scala 140:34:@1678.4]
  wire  _T_3506; // @[StoreQueue.scala 140:64:@1679.4]
  wire  _T_3510; // @[StoreQueue.scala 141:51:@1680.4]
  wire  _T_3511; // @[StoreQueue.scala 141:36:@1681.4]
  wire  noConflicts_15; // @[StoreQueue.scala 140:95:@1682.4]
  wire  _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_927; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _T_3519; // @[StoreQueue.scala 154:44:@1684.4]
  wire  _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _GEN_959; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3524; // @[StoreQueue.scala 154:66:@1685.4]
  wire  _T_3525; // @[StoreQueue.scala 154:63:@1686.4]
  wire  _T_3528; // @[StoreQueue.scala 154:109:@1688.4]
  wire  _T_3529; // @[StoreQueue.scala 154:109:@1689.4]
  wire  _T_3530; // @[StoreQueue.scala 154:109:@1690.4]
  wire  _T_3531; // @[StoreQueue.scala 154:109:@1691.4]
  wire  _T_3532; // @[StoreQueue.scala 154:109:@1692.4]
  wire  _T_3533; // @[StoreQueue.scala 154:109:@1693.4]
  wire  _T_3534; // @[StoreQueue.scala 154:109:@1694.4]
  wire  _T_3535; // @[StoreQueue.scala 154:109:@1695.4]
  wire  _T_3536; // @[StoreQueue.scala 154:109:@1696.4]
  wire  _T_3537; // @[StoreQueue.scala 154:109:@1697.4]
  wire  _T_3538; // @[StoreQueue.scala 154:109:@1698.4]
  wire  _T_3539; // @[StoreQueue.scala 154:109:@1699.4]
  wire  _T_3540; // @[StoreQueue.scala 154:109:@1700.4]
  wire  _T_3541; // @[StoreQueue.scala 154:109:@1701.4]
  wire  _T_3542; // @[StoreQueue.scala 154:109:@1702.4]
  wire  storeRequest; // @[StoreQueue.scala 154:88:@1703.4]
  wire  _T_3545; // @[StoreQueue.scala 164:23:@1708.6]
  wire  _T_3546; // @[StoreQueue.scala 164:43:@1709.6]
  wire  _T_3547; // @[StoreQueue.scala 164:59:@1710.6]
  wire  _GEN_960; // @[StoreQueue.scala 164:86:@1711.6]
  wire  _GEN_961; // @[StoreQueue.scala 162:37:@1704.4]
  wire  _T_3551; // @[StoreQueue.scala 164:23:@1718.6]
  wire  _T_3552; // @[StoreQueue.scala 164:43:@1719.6]
  wire  _T_3553; // @[StoreQueue.scala 164:59:@1720.6]
  wire  _GEN_962; // @[StoreQueue.scala 164:86:@1721.6]
  wire  _GEN_963; // @[StoreQueue.scala 162:37:@1714.4]
  wire  _T_3557; // @[StoreQueue.scala 164:23:@1728.6]
  wire  _T_3558; // @[StoreQueue.scala 164:43:@1729.6]
  wire  _T_3559; // @[StoreQueue.scala 164:59:@1730.6]
  wire  _GEN_964; // @[StoreQueue.scala 164:86:@1731.6]
  wire  _GEN_965; // @[StoreQueue.scala 162:37:@1724.4]
  wire  _T_3563; // @[StoreQueue.scala 164:23:@1738.6]
  wire  _T_3564; // @[StoreQueue.scala 164:43:@1739.6]
  wire  _T_3565; // @[StoreQueue.scala 164:59:@1740.6]
  wire  _GEN_966; // @[StoreQueue.scala 164:86:@1741.6]
  wire  _GEN_967; // @[StoreQueue.scala 162:37:@1734.4]
  wire  _T_3569; // @[StoreQueue.scala 164:23:@1748.6]
  wire  _T_3570; // @[StoreQueue.scala 164:43:@1749.6]
  wire  _T_3571; // @[StoreQueue.scala 164:59:@1750.6]
  wire  _GEN_968; // @[StoreQueue.scala 164:86:@1751.6]
  wire  _GEN_969; // @[StoreQueue.scala 162:37:@1744.4]
  wire  _T_3575; // @[StoreQueue.scala 164:23:@1758.6]
  wire  _T_3576; // @[StoreQueue.scala 164:43:@1759.6]
  wire  _T_3577; // @[StoreQueue.scala 164:59:@1760.6]
  wire  _GEN_970; // @[StoreQueue.scala 164:86:@1761.6]
  wire  _GEN_971; // @[StoreQueue.scala 162:37:@1754.4]
  wire  _T_3581; // @[StoreQueue.scala 164:23:@1768.6]
  wire  _T_3582; // @[StoreQueue.scala 164:43:@1769.6]
  wire  _T_3583; // @[StoreQueue.scala 164:59:@1770.6]
  wire  _GEN_972; // @[StoreQueue.scala 164:86:@1771.6]
  wire  _GEN_973; // @[StoreQueue.scala 162:37:@1764.4]
  wire  _T_3587; // @[StoreQueue.scala 164:23:@1778.6]
  wire  _T_3588; // @[StoreQueue.scala 164:43:@1779.6]
  wire  _T_3589; // @[StoreQueue.scala 164:59:@1780.6]
  wire  _GEN_974; // @[StoreQueue.scala 164:86:@1781.6]
  wire  _GEN_975; // @[StoreQueue.scala 162:37:@1774.4]
  wire  _T_3593; // @[StoreQueue.scala 164:23:@1788.6]
  wire  _T_3594; // @[StoreQueue.scala 164:43:@1789.6]
  wire  _T_3595; // @[StoreQueue.scala 164:59:@1790.6]
  wire  _GEN_976; // @[StoreQueue.scala 164:86:@1791.6]
  wire  _GEN_977; // @[StoreQueue.scala 162:37:@1784.4]
  wire  _T_3599; // @[StoreQueue.scala 164:23:@1798.6]
  wire  _T_3600; // @[StoreQueue.scala 164:43:@1799.6]
  wire  _T_3601; // @[StoreQueue.scala 164:59:@1800.6]
  wire  _GEN_978; // @[StoreQueue.scala 164:86:@1801.6]
  wire  _GEN_979; // @[StoreQueue.scala 162:37:@1794.4]
  wire  _T_3605; // @[StoreQueue.scala 164:23:@1808.6]
  wire  _T_3606; // @[StoreQueue.scala 164:43:@1809.6]
  wire  _T_3607; // @[StoreQueue.scala 164:59:@1810.6]
  wire  _GEN_980; // @[StoreQueue.scala 164:86:@1811.6]
  wire  _GEN_981; // @[StoreQueue.scala 162:37:@1804.4]
  wire  _T_3611; // @[StoreQueue.scala 164:23:@1818.6]
  wire  _T_3612; // @[StoreQueue.scala 164:43:@1819.6]
  wire  _T_3613; // @[StoreQueue.scala 164:59:@1820.6]
  wire  _GEN_982; // @[StoreQueue.scala 164:86:@1821.6]
  wire  _GEN_983; // @[StoreQueue.scala 162:37:@1814.4]
  wire  _T_3617; // @[StoreQueue.scala 164:23:@1828.6]
  wire  _T_3618; // @[StoreQueue.scala 164:43:@1829.6]
  wire  _T_3619; // @[StoreQueue.scala 164:59:@1830.6]
  wire  _GEN_984; // @[StoreQueue.scala 164:86:@1831.6]
  wire  _GEN_985; // @[StoreQueue.scala 162:37:@1824.4]
  wire  _T_3623; // @[StoreQueue.scala 164:23:@1838.6]
  wire  _T_3624; // @[StoreQueue.scala 164:43:@1839.6]
  wire  _T_3625; // @[StoreQueue.scala 164:59:@1840.6]
  wire  _GEN_986; // @[StoreQueue.scala 164:86:@1841.6]
  wire  _GEN_987; // @[StoreQueue.scala 162:37:@1834.4]
  wire  _T_3629; // @[StoreQueue.scala 164:23:@1848.6]
  wire  _T_3630; // @[StoreQueue.scala 164:43:@1849.6]
  wire  _T_3631; // @[StoreQueue.scala 164:59:@1850.6]
  wire  _GEN_988; // @[StoreQueue.scala 164:86:@1851.6]
  wire  _GEN_989; // @[StoreQueue.scala 162:37:@1844.4]
  wire  _T_3635; // @[StoreQueue.scala 164:23:@1858.6]
  wire  _T_3636; // @[StoreQueue.scala 164:43:@1859.6]
  wire  _T_3637; // @[StoreQueue.scala 164:59:@1860.6]
  wire  _GEN_990; // @[StoreQueue.scala 164:86:@1861.6]
  wire  _GEN_991; // @[StoreQueue.scala 162:37:@1854.4]
  wire  entriesPorts_0_0; // @[StoreQueue.scala 180:72:@1865.4]
  wire  entriesPorts_0_1; // @[StoreQueue.scala 180:72:@1867.4]
  wire  entriesPorts_0_2; // @[StoreQueue.scala 180:72:@1869.4]
  wire  entriesPorts_0_3; // @[StoreQueue.scala 180:72:@1871.4]
  wire  entriesPorts_0_4; // @[StoreQueue.scala 180:72:@1873.4]
  wire  entriesPorts_0_5; // @[StoreQueue.scala 180:72:@1875.4]
  wire  entriesPorts_0_6; // @[StoreQueue.scala 180:72:@1877.4]
  wire  entriesPorts_0_7; // @[StoreQueue.scala 180:72:@1879.4]
  wire  entriesPorts_0_8; // @[StoreQueue.scala 180:72:@1881.4]
  wire  entriesPorts_0_9; // @[StoreQueue.scala 180:72:@1883.4]
  wire  entriesPorts_0_10; // @[StoreQueue.scala 180:72:@1885.4]
  wire  entriesPorts_0_11; // @[StoreQueue.scala 180:72:@1887.4]
  wire  entriesPorts_0_12; // @[StoreQueue.scala 180:72:@1889.4]
  wire  entriesPorts_0_13; // @[StoreQueue.scala 180:72:@1891.4]
  wire  entriesPorts_0_14; // @[StoreQueue.scala 180:72:@1893.4]
  wire  entriesPorts_0_15; // @[StoreQueue.scala 180:72:@1895.4]
  wire  _T_4122; // @[StoreQueue.scala 192:91:@1899.4]
  wire  _T_4123; // @[StoreQueue.scala 192:88:@1900.4]
  wire  _T_4125; // @[StoreQueue.scala 192:91:@1901.4]
  wire  _T_4126; // @[StoreQueue.scala 192:88:@1902.4]
  wire  _T_4128; // @[StoreQueue.scala 192:91:@1903.4]
  wire  _T_4129; // @[StoreQueue.scala 192:88:@1904.4]
  wire  _T_4131; // @[StoreQueue.scala 192:91:@1905.4]
  wire  _T_4132; // @[StoreQueue.scala 192:88:@1906.4]
  wire  _T_4134; // @[StoreQueue.scala 192:91:@1907.4]
  wire  _T_4135; // @[StoreQueue.scala 192:88:@1908.4]
  wire  _T_4137; // @[StoreQueue.scala 192:91:@1909.4]
  wire  _T_4138; // @[StoreQueue.scala 192:88:@1910.4]
  wire  _T_4140; // @[StoreQueue.scala 192:91:@1911.4]
  wire  _T_4141; // @[StoreQueue.scala 192:88:@1912.4]
  wire  _T_4143; // @[StoreQueue.scala 192:91:@1913.4]
  wire  _T_4144; // @[StoreQueue.scala 192:88:@1914.4]
  wire  _T_4146; // @[StoreQueue.scala 192:91:@1915.4]
  wire  _T_4147; // @[StoreQueue.scala 192:88:@1916.4]
  wire  _T_4149; // @[StoreQueue.scala 192:91:@1917.4]
  wire  _T_4150; // @[StoreQueue.scala 192:88:@1918.4]
  wire  _T_4152; // @[StoreQueue.scala 192:91:@1919.4]
  wire  _T_4153; // @[StoreQueue.scala 192:88:@1920.4]
  wire  _T_4155; // @[StoreQueue.scala 192:91:@1921.4]
  wire  _T_4156; // @[StoreQueue.scala 192:88:@1922.4]
  wire  _T_4158; // @[StoreQueue.scala 192:91:@1923.4]
  wire  _T_4159; // @[StoreQueue.scala 192:88:@1924.4]
  wire  _T_4161; // @[StoreQueue.scala 192:91:@1925.4]
  wire  _T_4162; // @[StoreQueue.scala 192:88:@1926.4]
  wire  _T_4164; // @[StoreQueue.scala 192:91:@1927.4]
  wire  _T_4165; // @[StoreQueue.scala 192:88:@1928.4]
  wire  _T_4167; // @[StoreQueue.scala 192:91:@1929.4]
  wire  _T_4168; // @[StoreQueue.scala 192:88:@1930.4]
  wire  _T_4192; // @[StoreQueue.scala 193:91:@1948.4]
  wire  _T_4193; // @[StoreQueue.scala 193:88:@1949.4]
  wire  _T_4195; // @[StoreQueue.scala 193:91:@1950.4]
  wire  _T_4196; // @[StoreQueue.scala 193:88:@1951.4]
  wire  _T_4198; // @[StoreQueue.scala 193:91:@1952.4]
  wire  _T_4199; // @[StoreQueue.scala 193:88:@1953.4]
  wire  _T_4201; // @[StoreQueue.scala 193:91:@1954.4]
  wire  _T_4202; // @[StoreQueue.scala 193:88:@1955.4]
  wire  _T_4204; // @[StoreQueue.scala 193:91:@1956.4]
  wire  _T_4205; // @[StoreQueue.scala 193:88:@1957.4]
  wire  _T_4207; // @[StoreQueue.scala 193:91:@1958.4]
  wire  _T_4208; // @[StoreQueue.scala 193:88:@1959.4]
  wire  _T_4210; // @[StoreQueue.scala 193:91:@1960.4]
  wire  _T_4211; // @[StoreQueue.scala 193:88:@1961.4]
  wire  _T_4213; // @[StoreQueue.scala 193:91:@1962.4]
  wire  _T_4214; // @[StoreQueue.scala 193:88:@1963.4]
  wire  _T_4216; // @[StoreQueue.scala 193:91:@1964.4]
  wire  _T_4217; // @[StoreQueue.scala 193:88:@1965.4]
  wire  _T_4219; // @[StoreQueue.scala 193:91:@1966.4]
  wire  _T_4220; // @[StoreQueue.scala 193:88:@1967.4]
  wire  _T_4222; // @[StoreQueue.scala 193:91:@1968.4]
  wire  _T_4223; // @[StoreQueue.scala 193:88:@1969.4]
  wire  _T_4225; // @[StoreQueue.scala 193:91:@1970.4]
  wire  _T_4226; // @[StoreQueue.scala 193:88:@1971.4]
  wire  _T_4228; // @[StoreQueue.scala 193:91:@1972.4]
  wire  _T_4229; // @[StoreQueue.scala 193:88:@1973.4]
  wire  _T_4231; // @[StoreQueue.scala 193:91:@1974.4]
  wire  _T_4232; // @[StoreQueue.scala 193:88:@1975.4]
  wire  _T_4234; // @[StoreQueue.scala 193:91:@1976.4]
  wire  _T_4235; // @[StoreQueue.scala 193:88:@1977.4]
  wire  _T_4237; // @[StoreQueue.scala 193:91:@1978.4]
  wire  _T_4238; // @[StoreQueue.scala 193:88:@1979.4]
  wire [15:0] _T_4263; // @[OneHot.scala 52:12:@1998.4]
  wire  _T_4265; // @[util.scala 33:60:@2000.4]
  wire  _T_4266; // @[util.scala 33:60:@2001.4]
  wire  _T_4267; // @[util.scala 33:60:@2002.4]
  wire  _T_4268; // @[util.scala 33:60:@2003.4]
  wire  _T_4269; // @[util.scala 33:60:@2004.4]
  wire  _T_4270; // @[util.scala 33:60:@2005.4]
  wire  _T_4271; // @[util.scala 33:60:@2006.4]
  wire  _T_4272; // @[util.scala 33:60:@2007.4]
  wire  _T_4273; // @[util.scala 33:60:@2008.4]
  wire  _T_4274; // @[util.scala 33:60:@2009.4]
  wire  _T_4275; // @[util.scala 33:60:@2010.4]
  wire  _T_4276; // @[util.scala 33:60:@2011.4]
  wire  _T_4277; // @[util.scala 33:60:@2012.4]
  wire  _T_4278; // @[util.scala 33:60:@2013.4]
  wire  _T_4279; // @[util.scala 33:60:@2014.4]
  wire  _T_4280; // @[util.scala 33:60:@2015.4]
  wire [15:0] _T_4321; // @[Mux.scala 31:69:@2033.4]
  wire [15:0] _T_4322; // @[Mux.scala 31:69:@2034.4]
  wire [15:0] _T_4323; // @[Mux.scala 31:69:@2035.4]
  wire [15:0] _T_4324; // @[Mux.scala 31:69:@2036.4]
  wire [15:0] _T_4325; // @[Mux.scala 31:69:@2037.4]
  wire [15:0] _T_4326; // @[Mux.scala 31:69:@2038.4]
  wire [15:0] _T_4327; // @[Mux.scala 31:69:@2039.4]
  wire [15:0] _T_4328; // @[Mux.scala 31:69:@2040.4]
  wire [15:0] _T_4329; // @[Mux.scala 31:69:@2041.4]
  wire [15:0] _T_4330; // @[Mux.scala 31:69:@2042.4]
  wire [15:0] _T_4331; // @[Mux.scala 31:69:@2043.4]
  wire [15:0] _T_4332; // @[Mux.scala 31:69:@2044.4]
  wire [15:0] _T_4333; // @[Mux.scala 31:69:@2045.4]
  wire [15:0] _T_4334; // @[Mux.scala 31:69:@2046.4]
  wire [15:0] _T_4335; // @[Mux.scala 31:69:@2047.4]
  wire [15:0] _T_4336; // @[Mux.scala 31:69:@2048.4]
  wire  _T_4337; // @[OneHot.scala 66:30:@2049.4]
  wire  _T_4338; // @[OneHot.scala 66:30:@2050.4]
  wire  _T_4339; // @[OneHot.scala 66:30:@2051.4]
  wire  _T_4340; // @[OneHot.scala 66:30:@2052.4]
  wire  _T_4341; // @[OneHot.scala 66:30:@2053.4]
  wire  _T_4342; // @[OneHot.scala 66:30:@2054.4]
  wire  _T_4343; // @[OneHot.scala 66:30:@2055.4]
  wire  _T_4344; // @[OneHot.scala 66:30:@2056.4]
  wire  _T_4345; // @[OneHot.scala 66:30:@2057.4]
  wire  _T_4346; // @[OneHot.scala 66:30:@2058.4]
  wire  _T_4347; // @[OneHot.scala 66:30:@2059.4]
  wire  _T_4348; // @[OneHot.scala 66:30:@2060.4]
  wire  _T_4349; // @[OneHot.scala 66:30:@2061.4]
  wire  _T_4350; // @[OneHot.scala 66:30:@2062.4]
  wire  _T_4351; // @[OneHot.scala 66:30:@2063.4]
  wire  _T_4352; // @[OneHot.scala 66:30:@2064.4]
  wire [15:0] _T_4393; // @[Mux.scala 31:69:@2082.4]
  wire [15:0] _T_4394; // @[Mux.scala 31:69:@2083.4]
  wire [15:0] _T_4395; // @[Mux.scala 31:69:@2084.4]
  wire [15:0] _T_4396; // @[Mux.scala 31:69:@2085.4]
  wire [15:0] _T_4397; // @[Mux.scala 31:69:@2086.4]
  wire [15:0] _T_4398; // @[Mux.scala 31:69:@2087.4]
  wire [15:0] _T_4399; // @[Mux.scala 31:69:@2088.4]
  wire [15:0] _T_4400; // @[Mux.scala 31:69:@2089.4]
  wire [15:0] _T_4401; // @[Mux.scala 31:69:@2090.4]
  wire [15:0] _T_4402; // @[Mux.scala 31:69:@2091.4]
  wire [15:0] _T_4403; // @[Mux.scala 31:69:@2092.4]
  wire [15:0] _T_4404; // @[Mux.scala 31:69:@2093.4]
  wire [15:0] _T_4405; // @[Mux.scala 31:69:@2094.4]
  wire [15:0] _T_4406; // @[Mux.scala 31:69:@2095.4]
  wire [15:0] _T_4407; // @[Mux.scala 31:69:@2096.4]
  wire [15:0] _T_4408; // @[Mux.scala 31:69:@2097.4]
  wire  _T_4409; // @[OneHot.scala 66:30:@2098.4]
  wire  _T_4410; // @[OneHot.scala 66:30:@2099.4]
  wire  _T_4411; // @[OneHot.scala 66:30:@2100.4]
  wire  _T_4412; // @[OneHot.scala 66:30:@2101.4]
  wire  _T_4413; // @[OneHot.scala 66:30:@2102.4]
  wire  _T_4414; // @[OneHot.scala 66:30:@2103.4]
  wire  _T_4415; // @[OneHot.scala 66:30:@2104.4]
  wire  _T_4416; // @[OneHot.scala 66:30:@2105.4]
  wire  _T_4417; // @[OneHot.scala 66:30:@2106.4]
  wire  _T_4418; // @[OneHot.scala 66:30:@2107.4]
  wire  _T_4419; // @[OneHot.scala 66:30:@2108.4]
  wire  _T_4420; // @[OneHot.scala 66:30:@2109.4]
  wire  _T_4421; // @[OneHot.scala 66:30:@2110.4]
  wire  _T_4422; // @[OneHot.scala 66:30:@2111.4]
  wire  _T_4423; // @[OneHot.scala 66:30:@2112.4]
  wire  _T_4424; // @[OneHot.scala 66:30:@2113.4]
  wire [15:0] _T_4465; // @[Mux.scala 31:69:@2131.4]
  wire [15:0] _T_4466; // @[Mux.scala 31:69:@2132.4]
  wire [15:0] _T_4467; // @[Mux.scala 31:69:@2133.4]
  wire [15:0] _T_4468; // @[Mux.scala 31:69:@2134.4]
  wire [15:0] _T_4469; // @[Mux.scala 31:69:@2135.4]
  wire [15:0] _T_4470; // @[Mux.scala 31:69:@2136.4]
  wire [15:0] _T_4471; // @[Mux.scala 31:69:@2137.4]
  wire [15:0] _T_4472; // @[Mux.scala 31:69:@2138.4]
  wire [15:0] _T_4473; // @[Mux.scala 31:69:@2139.4]
  wire [15:0] _T_4474; // @[Mux.scala 31:69:@2140.4]
  wire [15:0] _T_4475; // @[Mux.scala 31:69:@2141.4]
  wire [15:0] _T_4476; // @[Mux.scala 31:69:@2142.4]
  wire [15:0] _T_4477; // @[Mux.scala 31:69:@2143.4]
  wire [15:0] _T_4478; // @[Mux.scala 31:69:@2144.4]
  wire [15:0] _T_4479; // @[Mux.scala 31:69:@2145.4]
  wire [15:0] _T_4480; // @[Mux.scala 31:69:@2146.4]
  wire  _T_4481; // @[OneHot.scala 66:30:@2147.4]
  wire  _T_4482; // @[OneHot.scala 66:30:@2148.4]
  wire  _T_4483; // @[OneHot.scala 66:30:@2149.4]
  wire  _T_4484; // @[OneHot.scala 66:30:@2150.4]
  wire  _T_4485; // @[OneHot.scala 66:30:@2151.4]
  wire  _T_4486; // @[OneHot.scala 66:30:@2152.4]
  wire  _T_4487; // @[OneHot.scala 66:30:@2153.4]
  wire  _T_4488; // @[OneHot.scala 66:30:@2154.4]
  wire  _T_4489; // @[OneHot.scala 66:30:@2155.4]
  wire  _T_4490; // @[OneHot.scala 66:30:@2156.4]
  wire  _T_4491; // @[OneHot.scala 66:30:@2157.4]
  wire  _T_4492; // @[OneHot.scala 66:30:@2158.4]
  wire  _T_4493; // @[OneHot.scala 66:30:@2159.4]
  wire  _T_4494; // @[OneHot.scala 66:30:@2160.4]
  wire  _T_4495; // @[OneHot.scala 66:30:@2161.4]
  wire  _T_4496; // @[OneHot.scala 66:30:@2162.4]
  wire [15:0] _T_4537; // @[Mux.scala 31:69:@2180.4]
  wire [15:0] _T_4538; // @[Mux.scala 31:69:@2181.4]
  wire [15:0] _T_4539; // @[Mux.scala 31:69:@2182.4]
  wire [15:0] _T_4540; // @[Mux.scala 31:69:@2183.4]
  wire [15:0] _T_4541; // @[Mux.scala 31:69:@2184.4]
  wire [15:0] _T_4542; // @[Mux.scala 31:69:@2185.4]
  wire [15:0] _T_4543; // @[Mux.scala 31:69:@2186.4]
  wire [15:0] _T_4544; // @[Mux.scala 31:69:@2187.4]
  wire [15:0] _T_4545; // @[Mux.scala 31:69:@2188.4]
  wire [15:0] _T_4546; // @[Mux.scala 31:69:@2189.4]
  wire [15:0] _T_4547; // @[Mux.scala 31:69:@2190.4]
  wire [15:0] _T_4548; // @[Mux.scala 31:69:@2191.4]
  wire [15:0] _T_4549; // @[Mux.scala 31:69:@2192.4]
  wire [15:0] _T_4550; // @[Mux.scala 31:69:@2193.4]
  wire [15:0] _T_4551; // @[Mux.scala 31:69:@2194.4]
  wire [15:0] _T_4552; // @[Mux.scala 31:69:@2195.4]
  wire  _T_4553; // @[OneHot.scala 66:30:@2196.4]
  wire  _T_4554; // @[OneHot.scala 66:30:@2197.4]
  wire  _T_4555; // @[OneHot.scala 66:30:@2198.4]
  wire  _T_4556; // @[OneHot.scala 66:30:@2199.4]
  wire  _T_4557; // @[OneHot.scala 66:30:@2200.4]
  wire  _T_4558; // @[OneHot.scala 66:30:@2201.4]
  wire  _T_4559; // @[OneHot.scala 66:30:@2202.4]
  wire  _T_4560; // @[OneHot.scala 66:30:@2203.4]
  wire  _T_4561; // @[OneHot.scala 66:30:@2204.4]
  wire  _T_4562; // @[OneHot.scala 66:30:@2205.4]
  wire  _T_4563; // @[OneHot.scala 66:30:@2206.4]
  wire  _T_4564; // @[OneHot.scala 66:30:@2207.4]
  wire  _T_4565; // @[OneHot.scala 66:30:@2208.4]
  wire  _T_4566; // @[OneHot.scala 66:30:@2209.4]
  wire  _T_4567; // @[OneHot.scala 66:30:@2210.4]
  wire  _T_4568; // @[OneHot.scala 66:30:@2211.4]
  wire [15:0] _T_4609; // @[Mux.scala 31:69:@2229.4]
  wire [15:0] _T_4610; // @[Mux.scala 31:69:@2230.4]
  wire [15:0] _T_4611; // @[Mux.scala 31:69:@2231.4]
  wire [15:0] _T_4612; // @[Mux.scala 31:69:@2232.4]
  wire [15:0] _T_4613; // @[Mux.scala 31:69:@2233.4]
  wire [15:0] _T_4614; // @[Mux.scala 31:69:@2234.4]
  wire [15:0] _T_4615; // @[Mux.scala 31:69:@2235.4]
  wire [15:0] _T_4616; // @[Mux.scala 31:69:@2236.4]
  wire [15:0] _T_4617; // @[Mux.scala 31:69:@2237.4]
  wire [15:0] _T_4618; // @[Mux.scala 31:69:@2238.4]
  wire [15:0] _T_4619; // @[Mux.scala 31:69:@2239.4]
  wire [15:0] _T_4620; // @[Mux.scala 31:69:@2240.4]
  wire [15:0] _T_4621; // @[Mux.scala 31:69:@2241.4]
  wire [15:0] _T_4622; // @[Mux.scala 31:69:@2242.4]
  wire [15:0] _T_4623; // @[Mux.scala 31:69:@2243.4]
  wire [15:0] _T_4624; // @[Mux.scala 31:69:@2244.4]
  wire  _T_4625; // @[OneHot.scala 66:30:@2245.4]
  wire  _T_4626; // @[OneHot.scala 66:30:@2246.4]
  wire  _T_4627; // @[OneHot.scala 66:30:@2247.4]
  wire  _T_4628; // @[OneHot.scala 66:30:@2248.4]
  wire  _T_4629; // @[OneHot.scala 66:30:@2249.4]
  wire  _T_4630; // @[OneHot.scala 66:30:@2250.4]
  wire  _T_4631; // @[OneHot.scala 66:30:@2251.4]
  wire  _T_4632; // @[OneHot.scala 66:30:@2252.4]
  wire  _T_4633; // @[OneHot.scala 66:30:@2253.4]
  wire  _T_4634; // @[OneHot.scala 66:30:@2254.4]
  wire  _T_4635; // @[OneHot.scala 66:30:@2255.4]
  wire  _T_4636; // @[OneHot.scala 66:30:@2256.4]
  wire  _T_4637; // @[OneHot.scala 66:30:@2257.4]
  wire  _T_4638; // @[OneHot.scala 66:30:@2258.4]
  wire  _T_4639; // @[OneHot.scala 66:30:@2259.4]
  wire  _T_4640; // @[OneHot.scala 66:30:@2260.4]
  wire [15:0] _T_4681; // @[Mux.scala 31:69:@2278.4]
  wire [15:0] _T_4682; // @[Mux.scala 31:69:@2279.4]
  wire [15:0] _T_4683; // @[Mux.scala 31:69:@2280.4]
  wire [15:0] _T_4684; // @[Mux.scala 31:69:@2281.4]
  wire [15:0] _T_4685; // @[Mux.scala 31:69:@2282.4]
  wire [15:0] _T_4686; // @[Mux.scala 31:69:@2283.4]
  wire [15:0] _T_4687; // @[Mux.scala 31:69:@2284.4]
  wire [15:0] _T_4688; // @[Mux.scala 31:69:@2285.4]
  wire [15:0] _T_4689; // @[Mux.scala 31:69:@2286.4]
  wire [15:0] _T_4690; // @[Mux.scala 31:69:@2287.4]
  wire [15:0] _T_4691; // @[Mux.scala 31:69:@2288.4]
  wire [15:0] _T_4692; // @[Mux.scala 31:69:@2289.4]
  wire [15:0] _T_4693; // @[Mux.scala 31:69:@2290.4]
  wire [15:0] _T_4694; // @[Mux.scala 31:69:@2291.4]
  wire [15:0] _T_4695; // @[Mux.scala 31:69:@2292.4]
  wire [15:0] _T_4696; // @[Mux.scala 31:69:@2293.4]
  wire  _T_4697; // @[OneHot.scala 66:30:@2294.4]
  wire  _T_4698; // @[OneHot.scala 66:30:@2295.4]
  wire  _T_4699; // @[OneHot.scala 66:30:@2296.4]
  wire  _T_4700; // @[OneHot.scala 66:30:@2297.4]
  wire  _T_4701; // @[OneHot.scala 66:30:@2298.4]
  wire  _T_4702; // @[OneHot.scala 66:30:@2299.4]
  wire  _T_4703; // @[OneHot.scala 66:30:@2300.4]
  wire  _T_4704; // @[OneHot.scala 66:30:@2301.4]
  wire  _T_4705; // @[OneHot.scala 66:30:@2302.4]
  wire  _T_4706; // @[OneHot.scala 66:30:@2303.4]
  wire  _T_4707; // @[OneHot.scala 66:30:@2304.4]
  wire  _T_4708; // @[OneHot.scala 66:30:@2305.4]
  wire  _T_4709; // @[OneHot.scala 66:30:@2306.4]
  wire  _T_4710; // @[OneHot.scala 66:30:@2307.4]
  wire  _T_4711; // @[OneHot.scala 66:30:@2308.4]
  wire  _T_4712; // @[OneHot.scala 66:30:@2309.4]
  wire [15:0] _T_4753; // @[Mux.scala 31:69:@2327.4]
  wire [15:0] _T_4754; // @[Mux.scala 31:69:@2328.4]
  wire [15:0] _T_4755; // @[Mux.scala 31:69:@2329.4]
  wire [15:0] _T_4756; // @[Mux.scala 31:69:@2330.4]
  wire [15:0] _T_4757; // @[Mux.scala 31:69:@2331.4]
  wire [15:0] _T_4758; // @[Mux.scala 31:69:@2332.4]
  wire [15:0] _T_4759; // @[Mux.scala 31:69:@2333.4]
  wire [15:0] _T_4760; // @[Mux.scala 31:69:@2334.4]
  wire [15:0] _T_4761; // @[Mux.scala 31:69:@2335.4]
  wire [15:0] _T_4762; // @[Mux.scala 31:69:@2336.4]
  wire [15:0] _T_4763; // @[Mux.scala 31:69:@2337.4]
  wire [15:0] _T_4764; // @[Mux.scala 31:69:@2338.4]
  wire [15:0] _T_4765; // @[Mux.scala 31:69:@2339.4]
  wire [15:0] _T_4766; // @[Mux.scala 31:69:@2340.4]
  wire [15:0] _T_4767; // @[Mux.scala 31:69:@2341.4]
  wire [15:0] _T_4768; // @[Mux.scala 31:69:@2342.4]
  wire  _T_4769; // @[OneHot.scala 66:30:@2343.4]
  wire  _T_4770; // @[OneHot.scala 66:30:@2344.4]
  wire  _T_4771; // @[OneHot.scala 66:30:@2345.4]
  wire  _T_4772; // @[OneHot.scala 66:30:@2346.4]
  wire  _T_4773; // @[OneHot.scala 66:30:@2347.4]
  wire  _T_4774; // @[OneHot.scala 66:30:@2348.4]
  wire  _T_4775; // @[OneHot.scala 66:30:@2349.4]
  wire  _T_4776; // @[OneHot.scala 66:30:@2350.4]
  wire  _T_4777; // @[OneHot.scala 66:30:@2351.4]
  wire  _T_4778; // @[OneHot.scala 66:30:@2352.4]
  wire  _T_4779; // @[OneHot.scala 66:30:@2353.4]
  wire  _T_4780; // @[OneHot.scala 66:30:@2354.4]
  wire  _T_4781; // @[OneHot.scala 66:30:@2355.4]
  wire  _T_4782; // @[OneHot.scala 66:30:@2356.4]
  wire  _T_4783; // @[OneHot.scala 66:30:@2357.4]
  wire  _T_4784; // @[OneHot.scala 66:30:@2358.4]
  wire [15:0] _T_4825; // @[Mux.scala 31:69:@2376.4]
  wire [15:0] _T_4826; // @[Mux.scala 31:69:@2377.4]
  wire [15:0] _T_4827; // @[Mux.scala 31:69:@2378.4]
  wire [15:0] _T_4828; // @[Mux.scala 31:69:@2379.4]
  wire [15:0] _T_4829; // @[Mux.scala 31:69:@2380.4]
  wire [15:0] _T_4830; // @[Mux.scala 31:69:@2381.4]
  wire [15:0] _T_4831; // @[Mux.scala 31:69:@2382.4]
  wire [15:0] _T_4832; // @[Mux.scala 31:69:@2383.4]
  wire [15:0] _T_4833; // @[Mux.scala 31:69:@2384.4]
  wire [15:0] _T_4834; // @[Mux.scala 31:69:@2385.4]
  wire [15:0] _T_4835; // @[Mux.scala 31:69:@2386.4]
  wire [15:0] _T_4836; // @[Mux.scala 31:69:@2387.4]
  wire [15:0] _T_4837; // @[Mux.scala 31:69:@2388.4]
  wire [15:0] _T_4838; // @[Mux.scala 31:69:@2389.4]
  wire [15:0] _T_4839; // @[Mux.scala 31:69:@2390.4]
  wire [15:0] _T_4840; // @[Mux.scala 31:69:@2391.4]
  wire  _T_4841; // @[OneHot.scala 66:30:@2392.4]
  wire  _T_4842; // @[OneHot.scala 66:30:@2393.4]
  wire  _T_4843; // @[OneHot.scala 66:30:@2394.4]
  wire  _T_4844; // @[OneHot.scala 66:30:@2395.4]
  wire  _T_4845; // @[OneHot.scala 66:30:@2396.4]
  wire  _T_4846; // @[OneHot.scala 66:30:@2397.4]
  wire  _T_4847; // @[OneHot.scala 66:30:@2398.4]
  wire  _T_4848; // @[OneHot.scala 66:30:@2399.4]
  wire  _T_4849; // @[OneHot.scala 66:30:@2400.4]
  wire  _T_4850; // @[OneHot.scala 66:30:@2401.4]
  wire  _T_4851; // @[OneHot.scala 66:30:@2402.4]
  wire  _T_4852; // @[OneHot.scala 66:30:@2403.4]
  wire  _T_4853; // @[OneHot.scala 66:30:@2404.4]
  wire  _T_4854; // @[OneHot.scala 66:30:@2405.4]
  wire  _T_4855; // @[OneHot.scala 66:30:@2406.4]
  wire  _T_4856; // @[OneHot.scala 66:30:@2407.4]
  wire [15:0] _T_4897; // @[Mux.scala 31:69:@2425.4]
  wire [15:0] _T_4898; // @[Mux.scala 31:69:@2426.4]
  wire [15:0] _T_4899; // @[Mux.scala 31:69:@2427.4]
  wire [15:0] _T_4900; // @[Mux.scala 31:69:@2428.4]
  wire [15:0] _T_4901; // @[Mux.scala 31:69:@2429.4]
  wire [15:0] _T_4902; // @[Mux.scala 31:69:@2430.4]
  wire [15:0] _T_4903; // @[Mux.scala 31:69:@2431.4]
  wire [15:0] _T_4904; // @[Mux.scala 31:69:@2432.4]
  wire [15:0] _T_4905; // @[Mux.scala 31:69:@2433.4]
  wire [15:0] _T_4906; // @[Mux.scala 31:69:@2434.4]
  wire [15:0] _T_4907; // @[Mux.scala 31:69:@2435.4]
  wire [15:0] _T_4908; // @[Mux.scala 31:69:@2436.4]
  wire [15:0] _T_4909; // @[Mux.scala 31:69:@2437.4]
  wire [15:0] _T_4910; // @[Mux.scala 31:69:@2438.4]
  wire [15:0] _T_4911; // @[Mux.scala 31:69:@2439.4]
  wire [15:0] _T_4912; // @[Mux.scala 31:69:@2440.4]
  wire  _T_4913; // @[OneHot.scala 66:30:@2441.4]
  wire  _T_4914; // @[OneHot.scala 66:30:@2442.4]
  wire  _T_4915; // @[OneHot.scala 66:30:@2443.4]
  wire  _T_4916; // @[OneHot.scala 66:30:@2444.4]
  wire  _T_4917; // @[OneHot.scala 66:30:@2445.4]
  wire  _T_4918; // @[OneHot.scala 66:30:@2446.4]
  wire  _T_4919; // @[OneHot.scala 66:30:@2447.4]
  wire  _T_4920; // @[OneHot.scala 66:30:@2448.4]
  wire  _T_4921; // @[OneHot.scala 66:30:@2449.4]
  wire  _T_4922; // @[OneHot.scala 66:30:@2450.4]
  wire  _T_4923; // @[OneHot.scala 66:30:@2451.4]
  wire  _T_4924; // @[OneHot.scala 66:30:@2452.4]
  wire  _T_4925; // @[OneHot.scala 66:30:@2453.4]
  wire  _T_4926; // @[OneHot.scala 66:30:@2454.4]
  wire  _T_4927; // @[OneHot.scala 66:30:@2455.4]
  wire  _T_4928; // @[OneHot.scala 66:30:@2456.4]
  wire [15:0] _T_4969; // @[Mux.scala 31:69:@2474.4]
  wire [15:0] _T_4970; // @[Mux.scala 31:69:@2475.4]
  wire [15:0] _T_4971; // @[Mux.scala 31:69:@2476.4]
  wire [15:0] _T_4972; // @[Mux.scala 31:69:@2477.4]
  wire [15:0] _T_4973; // @[Mux.scala 31:69:@2478.4]
  wire [15:0] _T_4974; // @[Mux.scala 31:69:@2479.4]
  wire [15:0] _T_4975; // @[Mux.scala 31:69:@2480.4]
  wire [15:0] _T_4976; // @[Mux.scala 31:69:@2481.4]
  wire [15:0] _T_4977; // @[Mux.scala 31:69:@2482.4]
  wire [15:0] _T_4978; // @[Mux.scala 31:69:@2483.4]
  wire [15:0] _T_4979; // @[Mux.scala 31:69:@2484.4]
  wire [15:0] _T_4980; // @[Mux.scala 31:69:@2485.4]
  wire [15:0] _T_4981; // @[Mux.scala 31:69:@2486.4]
  wire [15:0] _T_4982; // @[Mux.scala 31:69:@2487.4]
  wire [15:0] _T_4983; // @[Mux.scala 31:69:@2488.4]
  wire [15:0] _T_4984; // @[Mux.scala 31:69:@2489.4]
  wire  _T_4985; // @[OneHot.scala 66:30:@2490.4]
  wire  _T_4986; // @[OneHot.scala 66:30:@2491.4]
  wire  _T_4987; // @[OneHot.scala 66:30:@2492.4]
  wire  _T_4988; // @[OneHot.scala 66:30:@2493.4]
  wire  _T_4989; // @[OneHot.scala 66:30:@2494.4]
  wire  _T_4990; // @[OneHot.scala 66:30:@2495.4]
  wire  _T_4991; // @[OneHot.scala 66:30:@2496.4]
  wire  _T_4992; // @[OneHot.scala 66:30:@2497.4]
  wire  _T_4993; // @[OneHot.scala 66:30:@2498.4]
  wire  _T_4994; // @[OneHot.scala 66:30:@2499.4]
  wire  _T_4995; // @[OneHot.scala 66:30:@2500.4]
  wire  _T_4996; // @[OneHot.scala 66:30:@2501.4]
  wire  _T_4997; // @[OneHot.scala 66:30:@2502.4]
  wire  _T_4998; // @[OneHot.scala 66:30:@2503.4]
  wire  _T_4999; // @[OneHot.scala 66:30:@2504.4]
  wire  _T_5000; // @[OneHot.scala 66:30:@2505.4]
  wire [15:0] _T_5041; // @[Mux.scala 31:69:@2523.4]
  wire [15:0] _T_5042; // @[Mux.scala 31:69:@2524.4]
  wire [15:0] _T_5043; // @[Mux.scala 31:69:@2525.4]
  wire [15:0] _T_5044; // @[Mux.scala 31:69:@2526.4]
  wire [15:0] _T_5045; // @[Mux.scala 31:69:@2527.4]
  wire [15:0] _T_5046; // @[Mux.scala 31:69:@2528.4]
  wire [15:0] _T_5047; // @[Mux.scala 31:69:@2529.4]
  wire [15:0] _T_5048; // @[Mux.scala 31:69:@2530.4]
  wire [15:0] _T_5049; // @[Mux.scala 31:69:@2531.4]
  wire [15:0] _T_5050; // @[Mux.scala 31:69:@2532.4]
  wire [15:0] _T_5051; // @[Mux.scala 31:69:@2533.4]
  wire [15:0] _T_5052; // @[Mux.scala 31:69:@2534.4]
  wire [15:0] _T_5053; // @[Mux.scala 31:69:@2535.4]
  wire [15:0] _T_5054; // @[Mux.scala 31:69:@2536.4]
  wire [15:0] _T_5055; // @[Mux.scala 31:69:@2537.4]
  wire [15:0] _T_5056; // @[Mux.scala 31:69:@2538.4]
  wire  _T_5057; // @[OneHot.scala 66:30:@2539.4]
  wire  _T_5058; // @[OneHot.scala 66:30:@2540.4]
  wire  _T_5059; // @[OneHot.scala 66:30:@2541.4]
  wire  _T_5060; // @[OneHot.scala 66:30:@2542.4]
  wire  _T_5061; // @[OneHot.scala 66:30:@2543.4]
  wire  _T_5062; // @[OneHot.scala 66:30:@2544.4]
  wire  _T_5063; // @[OneHot.scala 66:30:@2545.4]
  wire  _T_5064; // @[OneHot.scala 66:30:@2546.4]
  wire  _T_5065; // @[OneHot.scala 66:30:@2547.4]
  wire  _T_5066; // @[OneHot.scala 66:30:@2548.4]
  wire  _T_5067; // @[OneHot.scala 66:30:@2549.4]
  wire  _T_5068; // @[OneHot.scala 66:30:@2550.4]
  wire  _T_5069; // @[OneHot.scala 66:30:@2551.4]
  wire  _T_5070; // @[OneHot.scala 66:30:@2552.4]
  wire  _T_5071; // @[OneHot.scala 66:30:@2553.4]
  wire  _T_5072; // @[OneHot.scala 66:30:@2554.4]
  wire [15:0] _T_5113; // @[Mux.scala 31:69:@2572.4]
  wire [15:0] _T_5114; // @[Mux.scala 31:69:@2573.4]
  wire [15:0] _T_5115; // @[Mux.scala 31:69:@2574.4]
  wire [15:0] _T_5116; // @[Mux.scala 31:69:@2575.4]
  wire [15:0] _T_5117; // @[Mux.scala 31:69:@2576.4]
  wire [15:0] _T_5118; // @[Mux.scala 31:69:@2577.4]
  wire [15:0] _T_5119; // @[Mux.scala 31:69:@2578.4]
  wire [15:0] _T_5120; // @[Mux.scala 31:69:@2579.4]
  wire [15:0] _T_5121; // @[Mux.scala 31:69:@2580.4]
  wire [15:0] _T_5122; // @[Mux.scala 31:69:@2581.4]
  wire [15:0] _T_5123; // @[Mux.scala 31:69:@2582.4]
  wire [15:0] _T_5124; // @[Mux.scala 31:69:@2583.4]
  wire [15:0] _T_5125; // @[Mux.scala 31:69:@2584.4]
  wire [15:0] _T_5126; // @[Mux.scala 31:69:@2585.4]
  wire [15:0] _T_5127; // @[Mux.scala 31:69:@2586.4]
  wire [15:0] _T_5128; // @[Mux.scala 31:69:@2587.4]
  wire  _T_5129; // @[OneHot.scala 66:30:@2588.4]
  wire  _T_5130; // @[OneHot.scala 66:30:@2589.4]
  wire  _T_5131; // @[OneHot.scala 66:30:@2590.4]
  wire  _T_5132; // @[OneHot.scala 66:30:@2591.4]
  wire  _T_5133; // @[OneHot.scala 66:30:@2592.4]
  wire  _T_5134; // @[OneHot.scala 66:30:@2593.4]
  wire  _T_5135; // @[OneHot.scala 66:30:@2594.4]
  wire  _T_5136; // @[OneHot.scala 66:30:@2595.4]
  wire  _T_5137; // @[OneHot.scala 66:30:@2596.4]
  wire  _T_5138; // @[OneHot.scala 66:30:@2597.4]
  wire  _T_5139; // @[OneHot.scala 66:30:@2598.4]
  wire  _T_5140; // @[OneHot.scala 66:30:@2599.4]
  wire  _T_5141; // @[OneHot.scala 66:30:@2600.4]
  wire  _T_5142; // @[OneHot.scala 66:30:@2601.4]
  wire  _T_5143; // @[OneHot.scala 66:30:@2602.4]
  wire  _T_5144; // @[OneHot.scala 66:30:@2603.4]
  wire [15:0] _T_5185; // @[Mux.scala 31:69:@2621.4]
  wire [15:0] _T_5186; // @[Mux.scala 31:69:@2622.4]
  wire [15:0] _T_5187; // @[Mux.scala 31:69:@2623.4]
  wire [15:0] _T_5188; // @[Mux.scala 31:69:@2624.4]
  wire [15:0] _T_5189; // @[Mux.scala 31:69:@2625.4]
  wire [15:0] _T_5190; // @[Mux.scala 31:69:@2626.4]
  wire [15:0] _T_5191; // @[Mux.scala 31:69:@2627.4]
  wire [15:0] _T_5192; // @[Mux.scala 31:69:@2628.4]
  wire [15:0] _T_5193; // @[Mux.scala 31:69:@2629.4]
  wire [15:0] _T_5194; // @[Mux.scala 31:69:@2630.4]
  wire [15:0] _T_5195; // @[Mux.scala 31:69:@2631.4]
  wire [15:0] _T_5196; // @[Mux.scala 31:69:@2632.4]
  wire [15:0] _T_5197; // @[Mux.scala 31:69:@2633.4]
  wire [15:0] _T_5198; // @[Mux.scala 31:69:@2634.4]
  wire [15:0] _T_5199; // @[Mux.scala 31:69:@2635.4]
  wire [15:0] _T_5200; // @[Mux.scala 31:69:@2636.4]
  wire  _T_5201; // @[OneHot.scala 66:30:@2637.4]
  wire  _T_5202; // @[OneHot.scala 66:30:@2638.4]
  wire  _T_5203; // @[OneHot.scala 66:30:@2639.4]
  wire  _T_5204; // @[OneHot.scala 66:30:@2640.4]
  wire  _T_5205; // @[OneHot.scala 66:30:@2641.4]
  wire  _T_5206; // @[OneHot.scala 66:30:@2642.4]
  wire  _T_5207; // @[OneHot.scala 66:30:@2643.4]
  wire  _T_5208; // @[OneHot.scala 66:30:@2644.4]
  wire  _T_5209; // @[OneHot.scala 66:30:@2645.4]
  wire  _T_5210; // @[OneHot.scala 66:30:@2646.4]
  wire  _T_5211; // @[OneHot.scala 66:30:@2647.4]
  wire  _T_5212; // @[OneHot.scala 66:30:@2648.4]
  wire  _T_5213; // @[OneHot.scala 66:30:@2649.4]
  wire  _T_5214; // @[OneHot.scala 66:30:@2650.4]
  wire  _T_5215; // @[OneHot.scala 66:30:@2651.4]
  wire  _T_5216; // @[OneHot.scala 66:30:@2652.4]
  wire [15:0] _T_5257; // @[Mux.scala 31:69:@2670.4]
  wire [15:0] _T_5258; // @[Mux.scala 31:69:@2671.4]
  wire [15:0] _T_5259; // @[Mux.scala 31:69:@2672.4]
  wire [15:0] _T_5260; // @[Mux.scala 31:69:@2673.4]
  wire [15:0] _T_5261; // @[Mux.scala 31:69:@2674.4]
  wire [15:0] _T_5262; // @[Mux.scala 31:69:@2675.4]
  wire [15:0] _T_5263; // @[Mux.scala 31:69:@2676.4]
  wire [15:0] _T_5264; // @[Mux.scala 31:69:@2677.4]
  wire [15:0] _T_5265; // @[Mux.scala 31:69:@2678.4]
  wire [15:0] _T_5266; // @[Mux.scala 31:69:@2679.4]
  wire [15:0] _T_5267; // @[Mux.scala 31:69:@2680.4]
  wire [15:0] _T_5268; // @[Mux.scala 31:69:@2681.4]
  wire [15:0] _T_5269; // @[Mux.scala 31:69:@2682.4]
  wire [15:0] _T_5270; // @[Mux.scala 31:69:@2683.4]
  wire [15:0] _T_5271; // @[Mux.scala 31:69:@2684.4]
  wire [15:0] _T_5272; // @[Mux.scala 31:69:@2685.4]
  wire  _T_5273; // @[OneHot.scala 66:30:@2686.4]
  wire  _T_5274; // @[OneHot.scala 66:30:@2687.4]
  wire  _T_5275; // @[OneHot.scala 66:30:@2688.4]
  wire  _T_5276; // @[OneHot.scala 66:30:@2689.4]
  wire  _T_5277; // @[OneHot.scala 66:30:@2690.4]
  wire  _T_5278; // @[OneHot.scala 66:30:@2691.4]
  wire  _T_5279; // @[OneHot.scala 66:30:@2692.4]
  wire  _T_5280; // @[OneHot.scala 66:30:@2693.4]
  wire  _T_5281; // @[OneHot.scala 66:30:@2694.4]
  wire  _T_5282; // @[OneHot.scala 66:30:@2695.4]
  wire  _T_5283; // @[OneHot.scala 66:30:@2696.4]
  wire  _T_5284; // @[OneHot.scala 66:30:@2697.4]
  wire  _T_5285; // @[OneHot.scala 66:30:@2698.4]
  wire  _T_5286; // @[OneHot.scala 66:30:@2699.4]
  wire  _T_5287; // @[OneHot.scala 66:30:@2700.4]
  wire  _T_5288; // @[OneHot.scala 66:30:@2701.4]
  wire [15:0] _T_5329; // @[Mux.scala 31:69:@2719.4]
  wire [15:0] _T_5330; // @[Mux.scala 31:69:@2720.4]
  wire [15:0] _T_5331; // @[Mux.scala 31:69:@2721.4]
  wire [15:0] _T_5332; // @[Mux.scala 31:69:@2722.4]
  wire [15:0] _T_5333; // @[Mux.scala 31:69:@2723.4]
  wire [15:0] _T_5334; // @[Mux.scala 31:69:@2724.4]
  wire [15:0] _T_5335; // @[Mux.scala 31:69:@2725.4]
  wire [15:0] _T_5336; // @[Mux.scala 31:69:@2726.4]
  wire [15:0] _T_5337; // @[Mux.scala 31:69:@2727.4]
  wire [15:0] _T_5338; // @[Mux.scala 31:69:@2728.4]
  wire [15:0] _T_5339; // @[Mux.scala 31:69:@2729.4]
  wire [15:0] _T_5340; // @[Mux.scala 31:69:@2730.4]
  wire [15:0] _T_5341; // @[Mux.scala 31:69:@2731.4]
  wire [15:0] _T_5342; // @[Mux.scala 31:69:@2732.4]
  wire [15:0] _T_5343; // @[Mux.scala 31:69:@2733.4]
  wire [15:0] _T_5344; // @[Mux.scala 31:69:@2734.4]
  wire  _T_5345; // @[OneHot.scala 66:30:@2735.4]
  wire  _T_5346; // @[OneHot.scala 66:30:@2736.4]
  wire  _T_5347; // @[OneHot.scala 66:30:@2737.4]
  wire  _T_5348; // @[OneHot.scala 66:30:@2738.4]
  wire  _T_5349; // @[OneHot.scala 66:30:@2739.4]
  wire  _T_5350; // @[OneHot.scala 66:30:@2740.4]
  wire  _T_5351; // @[OneHot.scala 66:30:@2741.4]
  wire  _T_5352; // @[OneHot.scala 66:30:@2742.4]
  wire  _T_5353; // @[OneHot.scala 66:30:@2743.4]
  wire  _T_5354; // @[OneHot.scala 66:30:@2744.4]
  wire  _T_5355; // @[OneHot.scala 66:30:@2745.4]
  wire  _T_5356; // @[OneHot.scala 66:30:@2746.4]
  wire  _T_5357; // @[OneHot.scala 66:30:@2747.4]
  wire  _T_5358; // @[OneHot.scala 66:30:@2748.4]
  wire  _T_5359; // @[OneHot.scala 66:30:@2749.4]
  wire  _T_5360; // @[OneHot.scala 66:30:@2750.4]
  wire [15:0] _T_5401; // @[Mux.scala 31:69:@2768.4]
  wire [15:0] _T_5402; // @[Mux.scala 31:69:@2769.4]
  wire [15:0] _T_5403; // @[Mux.scala 31:69:@2770.4]
  wire [15:0] _T_5404; // @[Mux.scala 31:69:@2771.4]
  wire [15:0] _T_5405; // @[Mux.scala 31:69:@2772.4]
  wire [15:0] _T_5406; // @[Mux.scala 31:69:@2773.4]
  wire [15:0] _T_5407; // @[Mux.scala 31:69:@2774.4]
  wire [15:0] _T_5408; // @[Mux.scala 31:69:@2775.4]
  wire [15:0] _T_5409; // @[Mux.scala 31:69:@2776.4]
  wire [15:0] _T_5410; // @[Mux.scala 31:69:@2777.4]
  wire [15:0] _T_5411; // @[Mux.scala 31:69:@2778.4]
  wire [15:0] _T_5412; // @[Mux.scala 31:69:@2779.4]
  wire [15:0] _T_5413; // @[Mux.scala 31:69:@2780.4]
  wire [15:0] _T_5414; // @[Mux.scala 31:69:@2781.4]
  wire [15:0] _T_5415; // @[Mux.scala 31:69:@2782.4]
  wire [15:0] _T_5416; // @[Mux.scala 31:69:@2783.4]
  wire  _T_5417; // @[OneHot.scala 66:30:@2784.4]
  wire  _T_5418; // @[OneHot.scala 66:30:@2785.4]
  wire  _T_5419; // @[OneHot.scala 66:30:@2786.4]
  wire  _T_5420; // @[OneHot.scala 66:30:@2787.4]
  wire  _T_5421; // @[OneHot.scala 66:30:@2788.4]
  wire  _T_5422; // @[OneHot.scala 66:30:@2789.4]
  wire  _T_5423; // @[OneHot.scala 66:30:@2790.4]
  wire  _T_5424; // @[OneHot.scala 66:30:@2791.4]
  wire  _T_5425; // @[OneHot.scala 66:30:@2792.4]
  wire  _T_5426; // @[OneHot.scala 66:30:@2793.4]
  wire  _T_5427; // @[OneHot.scala 66:30:@2794.4]
  wire  _T_5428; // @[OneHot.scala 66:30:@2795.4]
  wire  _T_5429; // @[OneHot.scala 66:30:@2796.4]
  wire  _T_5430; // @[OneHot.scala 66:30:@2797.4]
  wire  _T_5431; // @[OneHot.scala 66:30:@2798.4]
  wire  _T_5432; // @[OneHot.scala 66:30:@2799.4]
  wire [7:0] _T_5497; // @[Mux.scala 19:72:@2823.4]
  wire [15:0] _T_5505; // @[Mux.scala 19:72:@2831.4]
  wire [15:0] _T_5507; // @[Mux.scala 19:72:@2832.4]
  wire [7:0] _T_5514; // @[Mux.scala 19:72:@2839.4]
  wire [15:0] _T_5522; // @[Mux.scala 19:72:@2847.4]
  wire [15:0] _T_5524; // @[Mux.scala 19:72:@2848.4]
  wire [7:0] _T_5531; // @[Mux.scala 19:72:@2855.4]
  wire [15:0] _T_5539; // @[Mux.scala 19:72:@2863.4]
  wire [15:0] _T_5541; // @[Mux.scala 19:72:@2864.4]
  wire [7:0] _T_5548; // @[Mux.scala 19:72:@2871.4]
  wire [15:0] _T_5556; // @[Mux.scala 19:72:@2879.4]
  wire [15:0] _T_5558; // @[Mux.scala 19:72:@2880.4]
  wire [7:0] _T_5565; // @[Mux.scala 19:72:@2887.4]
  wire [15:0] _T_5573; // @[Mux.scala 19:72:@2895.4]
  wire [15:0] _T_5575; // @[Mux.scala 19:72:@2896.4]
  wire [7:0] _T_5582; // @[Mux.scala 19:72:@2903.4]
  wire [15:0] _T_5590; // @[Mux.scala 19:72:@2911.4]
  wire [15:0] _T_5592; // @[Mux.scala 19:72:@2912.4]
  wire [7:0] _T_5599; // @[Mux.scala 19:72:@2919.4]
  wire [15:0] _T_5607; // @[Mux.scala 19:72:@2927.4]
  wire [15:0] _T_5609; // @[Mux.scala 19:72:@2928.4]
  wire [7:0] _T_5616; // @[Mux.scala 19:72:@2935.4]
  wire [15:0] _T_5624; // @[Mux.scala 19:72:@2943.4]
  wire [15:0] _T_5626; // @[Mux.scala 19:72:@2944.4]
  wire [7:0] _T_5633; // @[Mux.scala 19:72:@2951.4]
  wire [15:0] _T_5641; // @[Mux.scala 19:72:@2959.4]
  wire [15:0] _T_5643; // @[Mux.scala 19:72:@2960.4]
  wire [7:0] _T_5650; // @[Mux.scala 19:72:@2967.4]
  wire [15:0] _T_5658; // @[Mux.scala 19:72:@2975.4]
  wire [15:0] _T_5660; // @[Mux.scala 19:72:@2976.4]
  wire [7:0] _T_5667; // @[Mux.scala 19:72:@2983.4]
  wire [15:0] _T_5675; // @[Mux.scala 19:72:@2991.4]
  wire [15:0] _T_5677; // @[Mux.scala 19:72:@2992.4]
  wire [7:0] _T_5684; // @[Mux.scala 19:72:@2999.4]
  wire [15:0] _T_5692; // @[Mux.scala 19:72:@3007.4]
  wire [15:0] _T_5694; // @[Mux.scala 19:72:@3008.4]
  wire [7:0] _T_5701; // @[Mux.scala 19:72:@3015.4]
  wire [15:0] _T_5709; // @[Mux.scala 19:72:@3023.4]
  wire [15:0] _T_5711; // @[Mux.scala 19:72:@3024.4]
  wire [7:0] _T_5718; // @[Mux.scala 19:72:@3031.4]
  wire [15:0] _T_5726; // @[Mux.scala 19:72:@3039.4]
  wire [15:0] _T_5728; // @[Mux.scala 19:72:@3040.4]
  wire [7:0] _T_5735; // @[Mux.scala 19:72:@3047.4]
  wire [15:0] _T_5743; // @[Mux.scala 19:72:@3055.4]
  wire [15:0] _T_5745; // @[Mux.scala 19:72:@3056.4]
  wire [7:0] _T_5752; // @[Mux.scala 19:72:@3063.4]
  wire [15:0] _T_5760; // @[Mux.scala 19:72:@3071.4]
  wire [15:0] _T_5762; // @[Mux.scala 19:72:@3072.4]
  wire [15:0] _T_5763; // @[Mux.scala 19:72:@3073.4]
  wire [15:0] _T_5764; // @[Mux.scala 19:72:@3074.4]
  wire [15:0] _T_5765; // @[Mux.scala 19:72:@3075.4]
  wire [15:0] _T_5766; // @[Mux.scala 19:72:@3076.4]
  wire [15:0] _T_5767; // @[Mux.scala 19:72:@3077.4]
  wire [15:0] _T_5768; // @[Mux.scala 19:72:@3078.4]
  wire [15:0] _T_5769; // @[Mux.scala 19:72:@3079.4]
  wire [15:0] _T_5770; // @[Mux.scala 19:72:@3080.4]
  wire [15:0] _T_5771; // @[Mux.scala 19:72:@3081.4]
  wire [15:0] _T_5772; // @[Mux.scala 19:72:@3082.4]
  wire [15:0] _T_5773; // @[Mux.scala 19:72:@3083.4]
  wire [15:0] _T_5774; // @[Mux.scala 19:72:@3084.4]
  wire [15:0] _T_5775; // @[Mux.scala 19:72:@3085.4]
  wire [15:0] _T_5776; // @[Mux.scala 19:72:@3086.4]
  wire [15:0] _T_5777; // @[Mux.scala 19:72:@3087.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@3091.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@3093.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@3095.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@3097.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@3099.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@3101.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@3103.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@3105.4]
  wire  inputAddrPriorityPorts_0_8; // @[Mux.scala 19:72:@3107.4]
  wire  inputAddrPriorityPorts_0_9; // @[Mux.scala 19:72:@3109.4]
  wire  inputAddrPriorityPorts_0_10; // @[Mux.scala 19:72:@3111.4]
  wire  inputAddrPriorityPorts_0_11; // @[Mux.scala 19:72:@3113.4]
  wire  inputAddrPriorityPorts_0_12; // @[Mux.scala 19:72:@3115.4]
  wire  inputAddrPriorityPorts_0_13; // @[Mux.scala 19:72:@3117.4]
  wire  inputAddrPriorityPorts_0_14; // @[Mux.scala 19:72:@3119.4]
  wire  inputAddrPriorityPorts_0_15; // @[Mux.scala 19:72:@3121.4]
  wire [15:0] _T_5979; // @[Mux.scala 31:69:@3175.4]
  wire [15:0] _T_5980; // @[Mux.scala 31:69:@3176.4]
  wire [15:0] _T_5981; // @[Mux.scala 31:69:@3177.4]
  wire [15:0] _T_5982; // @[Mux.scala 31:69:@3178.4]
  wire [15:0] _T_5983; // @[Mux.scala 31:69:@3179.4]
  wire [15:0] _T_5984; // @[Mux.scala 31:69:@3180.4]
  wire [15:0] _T_5985; // @[Mux.scala 31:69:@3181.4]
  wire [15:0] _T_5986; // @[Mux.scala 31:69:@3182.4]
  wire [15:0] _T_5987; // @[Mux.scala 31:69:@3183.4]
  wire [15:0] _T_5988; // @[Mux.scala 31:69:@3184.4]
  wire [15:0] _T_5989; // @[Mux.scala 31:69:@3185.4]
  wire [15:0] _T_5990; // @[Mux.scala 31:69:@3186.4]
  wire [15:0] _T_5991; // @[Mux.scala 31:69:@3187.4]
  wire [15:0] _T_5992; // @[Mux.scala 31:69:@3188.4]
  wire [15:0] _T_5993; // @[Mux.scala 31:69:@3189.4]
  wire [15:0] _T_5994; // @[Mux.scala 31:69:@3190.4]
  wire  _T_5995; // @[OneHot.scala 66:30:@3191.4]
  wire  _T_5996; // @[OneHot.scala 66:30:@3192.4]
  wire  _T_5997; // @[OneHot.scala 66:30:@3193.4]
  wire  _T_5998; // @[OneHot.scala 66:30:@3194.4]
  wire  _T_5999; // @[OneHot.scala 66:30:@3195.4]
  wire  _T_6000; // @[OneHot.scala 66:30:@3196.4]
  wire  _T_6001; // @[OneHot.scala 66:30:@3197.4]
  wire  _T_6002; // @[OneHot.scala 66:30:@3198.4]
  wire  _T_6003; // @[OneHot.scala 66:30:@3199.4]
  wire  _T_6004; // @[OneHot.scala 66:30:@3200.4]
  wire  _T_6005; // @[OneHot.scala 66:30:@3201.4]
  wire  _T_6006; // @[OneHot.scala 66:30:@3202.4]
  wire  _T_6007; // @[OneHot.scala 66:30:@3203.4]
  wire  _T_6008; // @[OneHot.scala 66:30:@3204.4]
  wire  _T_6009; // @[OneHot.scala 66:30:@3205.4]
  wire  _T_6010; // @[OneHot.scala 66:30:@3206.4]
  wire [15:0] _T_6051; // @[Mux.scala 31:69:@3224.4]
  wire [15:0] _T_6052; // @[Mux.scala 31:69:@3225.4]
  wire [15:0] _T_6053; // @[Mux.scala 31:69:@3226.4]
  wire [15:0] _T_6054; // @[Mux.scala 31:69:@3227.4]
  wire [15:0] _T_6055; // @[Mux.scala 31:69:@3228.4]
  wire [15:0] _T_6056; // @[Mux.scala 31:69:@3229.4]
  wire [15:0] _T_6057; // @[Mux.scala 31:69:@3230.4]
  wire [15:0] _T_6058; // @[Mux.scala 31:69:@3231.4]
  wire [15:0] _T_6059; // @[Mux.scala 31:69:@3232.4]
  wire [15:0] _T_6060; // @[Mux.scala 31:69:@3233.4]
  wire [15:0] _T_6061; // @[Mux.scala 31:69:@3234.4]
  wire [15:0] _T_6062; // @[Mux.scala 31:69:@3235.4]
  wire [15:0] _T_6063; // @[Mux.scala 31:69:@3236.4]
  wire [15:0] _T_6064; // @[Mux.scala 31:69:@3237.4]
  wire [15:0] _T_6065; // @[Mux.scala 31:69:@3238.4]
  wire [15:0] _T_6066; // @[Mux.scala 31:69:@3239.4]
  wire  _T_6067; // @[OneHot.scala 66:30:@3240.4]
  wire  _T_6068; // @[OneHot.scala 66:30:@3241.4]
  wire  _T_6069; // @[OneHot.scala 66:30:@3242.4]
  wire  _T_6070; // @[OneHot.scala 66:30:@3243.4]
  wire  _T_6071; // @[OneHot.scala 66:30:@3244.4]
  wire  _T_6072; // @[OneHot.scala 66:30:@3245.4]
  wire  _T_6073; // @[OneHot.scala 66:30:@3246.4]
  wire  _T_6074; // @[OneHot.scala 66:30:@3247.4]
  wire  _T_6075; // @[OneHot.scala 66:30:@3248.4]
  wire  _T_6076; // @[OneHot.scala 66:30:@3249.4]
  wire  _T_6077; // @[OneHot.scala 66:30:@3250.4]
  wire  _T_6078; // @[OneHot.scala 66:30:@3251.4]
  wire  _T_6079; // @[OneHot.scala 66:30:@3252.4]
  wire  _T_6080; // @[OneHot.scala 66:30:@3253.4]
  wire  _T_6081; // @[OneHot.scala 66:30:@3254.4]
  wire  _T_6082; // @[OneHot.scala 66:30:@3255.4]
  wire [15:0] _T_6123; // @[Mux.scala 31:69:@3273.4]
  wire [15:0] _T_6124; // @[Mux.scala 31:69:@3274.4]
  wire [15:0] _T_6125; // @[Mux.scala 31:69:@3275.4]
  wire [15:0] _T_6126; // @[Mux.scala 31:69:@3276.4]
  wire [15:0] _T_6127; // @[Mux.scala 31:69:@3277.4]
  wire [15:0] _T_6128; // @[Mux.scala 31:69:@3278.4]
  wire [15:0] _T_6129; // @[Mux.scala 31:69:@3279.4]
  wire [15:0] _T_6130; // @[Mux.scala 31:69:@3280.4]
  wire [15:0] _T_6131; // @[Mux.scala 31:69:@3281.4]
  wire [15:0] _T_6132; // @[Mux.scala 31:69:@3282.4]
  wire [15:0] _T_6133; // @[Mux.scala 31:69:@3283.4]
  wire [15:0] _T_6134; // @[Mux.scala 31:69:@3284.4]
  wire [15:0] _T_6135; // @[Mux.scala 31:69:@3285.4]
  wire [15:0] _T_6136; // @[Mux.scala 31:69:@3286.4]
  wire [15:0] _T_6137; // @[Mux.scala 31:69:@3287.4]
  wire [15:0] _T_6138; // @[Mux.scala 31:69:@3288.4]
  wire  _T_6139; // @[OneHot.scala 66:30:@3289.4]
  wire  _T_6140; // @[OneHot.scala 66:30:@3290.4]
  wire  _T_6141; // @[OneHot.scala 66:30:@3291.4]
  wire  _T_6142; // @[OneHot.scala 66:30:@3292.4]
  wire  _T_6143; // @[OneHot.scala 66:30:@3293.4]
  wire  _T_6144; // @[OneHot.scala 66:30:@3294.4]
  wire  _T_6145; // @[OneHot.scala 66:30:@3295.4]
  wire  _T_6146; // @[OneHot.scala 66:30:@3296.4]
  wire  _T_6147; // @[OneHot.scala 66:30:@3297.4]
  wire  _T_6148; // @[OneHot.scala 66:30:@3298.4]
  wire  _T_6149; // @[OneHot.scala 66:30:@3299.4]
  wire  _T_6150; // @[OneHot.scala 66:30:@3300.4]
  wire  _T_6151; // @[OneHot.scala 66:30:@3301.4]
  wire  _T_6152; // @[OneHot.scala 66:30:@3302.4]
  wire  _T_6153; // @[OneHot.scala 66:30:@3303.4]
  wire  _T_6154; // @[OneHot.scala 66:30:@3304.4]
  wire [15:0] _T_6195; // @[Mux.scala 31:69:@3322.4]
  wire [15:0] _T_6196; // @[Mux.scala 31:69:@3323.4]
  wire [15:0] _T_6197; // @[Mux.scala 31:69:@3324.4]
  wire [15:0] _T_6198; // @[Mux.scala 31:69:@3325.4]
  wire [15:0] _T_6199; // @[Mux.scala 31:69:@3326.4]
  wire [15:0] _T_6200; // @[Mux.scala 31:69:@3327.4]
  wire [15:0] _T_6201; // @[Mux.scala 31:69:@3328.4]
  wire [15:0] _T_6202; // @[Mux.scala 31:69:@3329.4]
  wire [15:0] _T_6203; // @[Mux.scala 31:69:@3330.4]
  wire [15:0] _T_6204; // @[Mux.scala 31:69:@3331.4]
  wire [15:0] _T_6205; // @[Mux.scala 31:69:@3332.4]
  wire [15:0] _T_6206; // @[Mux.scala 31:69:@3333.4]
  wire [15:0] _T_6207; // @[Mux.scala 31:69:@3334.4]
  wire [15:0] _T_6208; // @[Mux.scala 31:69:@3335.4]
  wire [15:0] _T_6209; // @[Mux.scala 31:69:@3336.4]
  wire [15:0] _T_6210; // @[Mux.scala 31:69:@3337.4]
  wire  _T_6211; // @[OneHot.scala 66:30:@3338.4]
  wire  _T_6212; // @[OneHot.scala 66:30:@3339.4]
  wire  _T_6213; // @[OneHot.scala 66:30:@3340.4]
  wire  _T_6214; // @[OneHot.scala 66:30:@3341.4]
  wire  _T_6215; // @[OneHot.scala 66:30:@3342.4]
  wire  _T_6216; // @[OneHot.scala 66:30:@3343.4]
  wire  _T_6217; // @[OneHot.scala 66:30:@3344.4]
  wire  _T_6218; // @[OneHot.scala 66:30:@3345.4]
  wire  _T_6219; // @[OneHot.scala 66:30:@3346.4]
  wire  _T_6220; // @[OneHot.scala 66:30:@3347.4]
  wire  _T_6221; // @[OneHot.scala 66:30:@3348.4]
  wire  _T_6222; // @[OneHot.scala 66:30:@3349.4]
  wire  _T_6223; // @[OneHot.scala 66:30:@3350.4]
  wire  _T_6224; // @[OneHot.scala 66:30:@3351.4]
  wire  _T_6225; // @[OneHot.scala 66:30:@3352.4]
  wire  _T_6226; // @[OneHot.scala 66:30:@3353.4]
  wire [15:0] _T_6267; // @[Mux.scala 31:69:@3371.4]
  wire [15:0] _T_6268; // @[Mux.scala 31:69:@3372.4]
  wire [15:0] _T_6269; // @[Mux.scala 31:69:@3373.4]
  wire [15:0] _T_6270; // @[Mux.scala 31:69:@3374.4]
  wire [15:0] _T_6271; // @[Mux.scala 31:69:@3375.4]
  wire [15:0] _T_6272; // @[Mux.scala 31:69:@3376.4]
  wire [15:0] _T_6273; // @[Mux.scala 31:69:@3377.4]
  wire [15:0] _T_6274; // @[Mux.scala 31:69:@3378.4]
  wire [15:0] _T_6275; // @[Mux.scala 31:69:@3379.4]
  wire [15:0] _T_6276; // @[Mux.scala 31:69:@3380.4]
  wire [15:0] _T_6277; // @[Mux.scala 31:69:@3381.4]
  wire [15:0] _T_6278; // @[Mux.scala 31:69:@3382.4]
  wire [15:0] _T_6279; // @[Mux.scala 31:69:@3383.4]
  wire [15:0] _T_6280; // @[Mux.scala 31:69:@3384.4]
  wire [15:0] _T_6281; // @[Mux.scala 31:69:@3385.4]
  wire [15:0] _T_6282; // @[Mux.scala 31:69:@3386.4]
  wire  _T_6283; // @[OneHot.scala 66:30:@3387.4]
  wire  _T_6284; // @[OneHot.scala 66:30:@3388.4]
  wire  _T_6285; // @[OneHot.scala 66:30:@3389.4]
  wire  _T_6286; // @[OneHot.scala 66:30:@3390.4]
  wire  _T_6287; // @[OneHot.scala 66:30:@3391.4]
  wire  _T_6288; // @[OneHot.scala 66:30:@3392.4]
  wire  _T_6289; // @[OneHot.scala 66:30:@3393.4]
  wire  _T_6290; // @[OneHot.scala 66:30:@3394.4]
  wire  _T_6291; // @[OneHot.scala 66:30:@3395.4]
  wire  _T_6292; // @[OneHot.scala 66:30:@3396.4]
  wire  _T_6293; // @[OneHot.scala 66:30:@3397.4]
  wire  _T_6294; // @[OneHot.scala 66:30:@3398.4]
  wire  _T_6295; // @[OneHot.scala 66:30:@3399.4]
  wire  _T_6296; // @[OneHot.scala 66:30:@3400.4]
  wire  _T_6297; // @[OneHot.scala 66:30:@3401.4]
  wire  _T_6298; // @[OneHot.scala 66:30:@3402.4]
  wire [15:0] _T_6339; // @[Mux.scala 31:69:@3420.4]
  wire [15:0] _T_6340; // @[Mux.scala 31:69:@3421.4]
  wire [15:0] _T_6341; // @[Mux.scala 31:69:@3422.4]
  wire [15:0] _T_6342; // @[Mux.scala 31:69:@3423.4]
  wire [15:0] _T_6343; // @[Mux.scala 31:69:@3424.4]
  wire [15:0] _T_6344; // @[Mux.scala 31:69:@3425.4]
  wire [15:0] _T_6345; // @[Mux.scala 31:69:@3426.4]
  wire [15:0] _T_6346; // @[Mux.scala 31:69:@3427.4]
  wire [15:0] _T_6347; // @[Mux.scala 31:69:@3428.4]
  wire [15:0] _T_6348; // @[Mux.scala 31:69:@3429.4]
  wire [15:0] _T_6349; // @[Mux.scala 31:69:@3430.4]
  wire [15:0] _T_6350; // @[Mux.scala 31:69:@3431.4]
  wire [15:0] _T_6351; // @[Mux.scala 31:69:@3432.4]
  wire [15:0] _T_6352; // @[Mux.scala 31:69:@3433.4]
  wire [15:0] _T_6353; // @[Mux.scala 31:69:@3434.4]
  wire [15:0] _T_6354; // @[Mux.scala 31:69:@3435.4]
  wire  _T_6355; // @[OneHot.scala 66:30:@3436.4]
  wire  _T_6356; // @[OneHot.scala 66:30:@3437.4]
  wire  _T_6357; // @[OneHot.scala 66:30:@3438.4]
  wire  _T_6358; // @[OneHot.scala 66:30:@3439.4]
  wire  _T_6359; // @[OneHot.scala 66:30:@3440.4]
  wire  _T_6360; // @[OneHot.scala 66:30:@3441.4]
  wire  _T_6361; // @[OneHot.scala 66:30:@3442.4]
  wire  _T_6362; // @[OneHot.scala 66:30:@3443.4]
  wire  _T_6363; // @[OneHot.scala 66:30:@3444.4]
  wire  _T_6364; // @[OneHot.scala 66:30:@3445.4]
  wire  _T_6365; // @[OneHot.scala 66:30:@3446.4]
  wire  _T_6366; // @[OneHot.scala 66:30:@3447.4]
  wire  _T_6367; // @[OneHot.scala 66:30:@3448.4]
  wire  _T_6368; // @[OneHot.scala 66:30:@3449.4]
  wire  _T_6369; // @[OneHot.scala 66:30:@3450.4]
  wire  _T_6370; // @[OneHot.scala 66:30:@3451.4]
  wire [15:0] _T_6411; // @[Mux.scala 31:69:@3469.4]
  wire [15:0] _T_6412; // @[Mux.scala 31:69:@3470.4]
  wire [15:0] _T_6413; // @[Mux.scala 31:69:@3471.4]
  wire [15:0] _T_6414; // @[Mux.scala 31:69:@3472.4]
  wire [15:0] _T_6415; // @[Mux.scala 31:69:@3473.4]
  wire [15:0] _T_6416; // @[Mux.scala 31:69:@3474.4]
  wire [15:0] _T_6417; // @[Mux.scala 31:69:@3475.4]
  wire [15:0] _T_6418; // @[Mux.scala 31:69:@3476.4]
  wire [15:0] _T_6419; // @[Mux.scala 31:69:@3477.4]
  wire [15:0] _T_6420; // @[Mux.scala 31:69:@3478.4]
  wire [15:0] _T_6421; // @[Mux.scala 31:69:@3479.4]
  wire [15:0] _T_6422; // @[Mux.scala 31:69:@3480.4]
  wire [15:0] _T_6423; // @[Mux.scala 31:69:@3481.4]
  wire [15:0] _T_6424; // @[Mux.scala 31:69:@3482.4]
  wire [15:0] _T_6425; // @[Mux.scala 31:69:@3483.4]
  wire [15:0] _T_6426; // @[Mux.scala 31:69:@3484.4]
  wire  _T_6427; // @[OneHot.scala 66:30:@3485.4]
  wire  _T_6428; // @[OneHot.scala 66:30:@3486.4]
  wire  _T_6429; // @[OneHot.scala 66:30:@3487.4]
  wire  _T_6430; // @[OneHot.scala 66:30:@3488.4]
  wire  _T_6431; // @[OneHot.scala 66:30:@3489.4]
  wire  _T_6432; // @[OneHot.scala 66:30:@3490.4]
  wire  _T_6433; // @[OneHot.scala 66:30:@3491.4]
  wire  _T_6434; // @[OneHot.scala 66:30:@3492.4]
  wire  _T_6435; // @[OneHot.scala 66:30:@3493.4]
  wire  _T_6436; // @[OneHot.scala 66:30:@3494.4]
  wire  _T_6437; // @[OneHot.scala 66:30:@3495.4]
  wire  _T_6438; // @[OneHot.scala 66:30:@3496.4]
  wire  _T_6439; // @[OneHot.scala 66:30:@3497.4]
  wire  _T_6440; // @[OneHot.scala 66:30:@3498.4]
  wire  _T_6441; // @[OneHot.scala 66:30:@3499.4]
  wire  _T_6442; // @[OneHot.scala 66:30:@3500.4]
  wire [15:0] _T_6483; // @[Mux.scala 31:69:@3518.4]
  wire [15:0] _T_6484; // @[Mux.scala 31:69:@3519.4]
  wire [15:0] _T_6485; // @[Mux.scala 31:69:@3520.4]
  wire [15:0] _T_6486; // @[Mux.scala 31:69:@3521.4]
  wire [15:0] _T_6487; // @[Mux.scala 31:69:@3522.4]
  wire [15:0] _T_6488; // @[Mux.scala 31:69:@3523.4]
  wire [15:0] _T_6489; // @[Mux.scala 31:69:@3524.4]
  wire [15:0] _T_6490; // @[Mux.scala 31:69:@3525.4]
  wire [15:0] _T_6491; // @[Mux.scala 31:69:@3526.4]
  wire [15:0] _T_6492; // @[Mux.scala 31:69:@3527.4]
  wire [15:0] _T_6493; // @[Mux.scala 31:69:@3528.4]
  wire [15:0] _T_6494; // @[Mux.scala 31:69:@3529.4]
  wire [15:0] _T_6495; // @[Mux.scala 31:69:@3530.4]
  wire [15:0] _T_6496; // @[Mux.scala 31:69:@3531.4]
  wire [15:0] _T_6497; // @[Mux.scala 31:69:@3532.4]
  wire [15:0] _T_6498; // @[Mux.scala 31:69:@3533.4]
  wire  _T_6499; // @[OneHot.scala 66:30:@3534.4]
  wire  _T_6500; // @[OneHot.scala 66:30:@3535.4]
  wire  _T_6501; // @[OneHot.scala 66:30:@3536.4]
  wire  _T_6502; // @[OneHot.scala 66:30:@3537.4]
  wire  _T_6503; // @[OneHot.scala 66:30:@3538.4]
  wire  _T_6504; // @[OneHot.scala 66:30:@3539.4]
  wire  _T_6505; // @[OneHot.scala 66:30:@3540.4]
  wire  _T_6506; // @[OneHot.scala 66:30:@3541.4]
  wire  _T_6507; // @[OneHot.scala 66:30:@3542.4]
  wire  _T_6508; // @[OneHot.scala 66:30:@3543.4]
  wire  _T_6509; // @[OneHot.scala 66:30:@3544.4]
  wire  _T_6510; // @[OneHot.scala 66:30:@3545.4]
  wire  _T_6511; // @[OneHot.scala 66:30:@3546.4]
  wire  _T_6512; // @[OneHot.scala 66:30:@3547.4]
  wire  _T_6513; // @[OneHot.scala 66:30:@3548.4]
  wire  _T_6514; // @[OneHot.scala 66:30:@3549.4]
  wire [15:0] _T_6555; // @[Mux.scala 31:69:@3567.4]
  wire [15:0] _T_6556; // @[Mux.scala 31:69:@3568.4]
  wire [15:0] _T_6557; // @[Mux.scala 31:69:@3569.4]
  wire [15:0] _T_6558; // @[Mux.scala 31:69:@3570.4]
  wire [15:0] _T_6559; // @[Mux.scala 31:69:@3571.4]
  wire [15:0] _T_6560; // @[Mux.scala 31:69:@3572.4]
  wire [15:0] _T_6561; // @[Mux.scala 31:69:@3573.4]
  wire [15:0] _T_6562; // @[Mux.scala 31:69:@3574.4]
  wire [15:0] _T_6563; // @[Mux.scala 31:69:@3575.4]
  wire [15:0] _T_6564; // @[Mux.scala 31:69:@3576.4]
  wire [15:0] _T_6565; // @[Mux.scala 31:69:@3577.4]
  wire [15:0] _T_6566; // @[Mux.scala 31:69:@3578.4]
  wire [15:0] _T_6567; // @[Mux.scala 31:69:@3579.4]
  wire [15:0] _T_6568; // @[Mux.scala 31:69:@3580.4]
  wire [15:0] _T_6569; // @[Mux.scala 31:69:@3581.4]
  wire [15:0] _T_6570; // @[Mux.scala 31:69:@3582.4]
  wire  _T_6571; // @[OneHot.scala 66:30:@3583.4]
  wire  _T_6572; // @[OneHot.scala 66:30:@3584.4]
  wire  _T_6573; // @[OneHot.scala 66:30:@3585.4]
  wire  _T_6574; // @[OneHot.scala 66:30:@3586.4]
  wire  _T_6575; // @[OneHot.scala 66:30:@3587.4]
  wire  _T_6576; // @[OneHot.scala 66:30:@3588.4]
  wire  _T_6577; // @[OneHot.scala 66:30:@3589.4]
  wire  _T_6578; // @[OneHot.scala 66:30:@3590.4]
  wire  _T_6579; // @[OneHot.scala 66:30:@3591.4]
  wire  _T_6580; // @[OneHot.scala 66:30:@3592.4]
  wire  _T_6581; // @[OneHot.scala 66:30:@3593.4]
  wire  _T_6582; // @[OneHot.scala 66:30:@3594.4]
  wire  _T_6583; // @[OneHot.scala 66:30:@3595.4]
  wire  _T_6584; // @[OneHot.scala 66:30:@3596.4]
  wire  _T_6585; // @[OneHot.scala 66:30:@3597.4]
  wire  _T_6586; // @[OneHot.scala 66:30:@3598.4]
  wire [15:0] _T_6627; // @[Mux.scala 31:69:@3616.4]
  wire [15:0] _T_6628; // @[Mux.scala 31:69:@3617.4]
  wire [15:0] _T_6629; // @[Mux.scala 31:69:@3618.4]
  wire [15:0] _T_6630; // @[Mux.scala 31:69:@3619.4]
  wire [15:0] _T_6631; // @[Mux.scala 31:69:@3620.4]
  wire [15:0] _T_6632; // @[Mux.scala 31:69:@3621.4]
  wire [15:0] _T_6633; // @[Mux.scala 31:69:@3622.4]
  wire [15:0] _T_6634; // @[Mux.scala 31:69:@3623.4]
  wire [15:0] _T_6635; // @[Mux.scala 31:69:@3624.4]
  wire [15:0] _T_6636; // @[Mux.scala 31:69:@3625.4]
  wire [15:0] _T_6637; // @[Mux.scala 31:69:@3626.4]
  wire [15:0] _T_6638; // @[Mux.scala 31:69:@3627.4]
  wire [15:0] _T_6639; // @[Mux.scala 31:69:@3628.4]
  wire [15:0] _T_6640; // @[Mux.scala 31:69:@3629.4]
  wire [15:0] _T_6641; // @[Mux.scala 31:69:@3630.4]
  wire [15:0] _T_6642; // @[Mux.scala 31:69:@3631.4]
  wire  _T_6643; // @[OneHot.scala 66:30:@3632.4]
  wire  _T_6644; // @[OneHot.scala 66:30:@3633.4]
  wire  _T_6645; // @[OneHot.scala 66:30:@3634.4]
  wire  _T_6646; // @[OneHot.scala 66:30:@3635.4]
  wire  _T_6647; // @[OneHot.scala 66:30:@3636.4]
  wire  _T_6648; // @[OneHot.scala 66:30:@3637.4]
  wire  _T_6649; // @[OneHot.scala 66:30:@3638.4]
  wire  _T_6650; // @[OneHot.scala 66:30:@3639.4]
  wire  _T_6651; // @[OneHot.scala 66:30:@3640.4]
  wire  _T_6652; // @[OneHot.scala 66:30:@3641.4]
  wire  _T_6653; // @[OneHot.scala 66:30:@3642.4]
  wire  _T_6654; // @[OneHot.scala 66:30:@3643.4]
  wire  _T_6655; // @[OneHot.scala 66:30:@3644.4]
  wire  _T_6656; // @[OneHot.scala 66:30:@3645.4]
  wire  _T_6657; // @[OneHot.scala 66:30:@3646.4]
  wire  _T_6658; // @[OneHot.scala 66:30:@3647.4]
  wire [15:0] _T_6699; // @[Mux.scala 31:69:@3665.4]
  wire [15:0] _T_6700; // @[Mux.scala 31:69:@3666.4]
  wire [15:0] _T_6701; // @[Mux.scala 31:69:@3667.4]
  wire [15:0] _T_6702; // @[Mux.scala 31:69:@3668.4]
  wire [15:0] _T_6703; // @[Mux.scala 31:69:@3669.4]
  wire [15:0] _T_6704; // @[Mux.scala 31:69:@3670.4]
  wire [15:0] _T_6705; // @[Mux.scala 31:69:@3671.4]
  wire [15:0] _T_6706; // @[Mux.scala 31:69:@3672.4]
  wire [15:0] _T_6707; // @[Mux.scala 31:69:@3673.4]
  wire [15:0] _T_6708; // @[Mux.scala 31:69:@3674.4]
  wire [15:0] _T_6709; // @[Mux.scala 31:69:@3675.4]
  wire [15:0] _T_6710; // @[Mux.scala 31:69:@3676.4]
  wire [15:0] _T_6711; // @[Mux.scala 31:69:@3677.4]
  wire [15:0] _T_6712; // @[Mux.scala 31:69:@3678.4]
  wire [15:0] _T_6713; // @[Mux.scala 31:69:@3679.4]
  wire [15:0] _T_6714; // @[Mux.scala 31:69:@3680.4]
  wire  _T_6715; // @[OneHot.scala 66:30:@3681.4]
  wire  _T_6716; // @[OneHot.scala 66:30:@3682.4]
  wire  _T_6717; // @[OneHot.scala 66:30:@3683.4]
  wire  _T_6718; // @[OneHot.scala 66:30:@3684.4]
  wire  _T_6719; // @[OneHot.scala 66:30:@3685.4]
  wire  _T_6720; // @[OneHot.scala 66:30:@3686.4]
  wire  _T_6721; // @[OneHot.scala 66:30:@3687.4]
  wire  _T_6722; // @[OneHot.scala 66:30:@3688.4]
  wire  _T_6723; // @[OneHot.scala 66:30:@3689.4]
  wire  _T_6724; // @[OneHot.scala 66:30:@3690.4]
  wire  _T_6725; // @[OneHot.scala 66:30:@3691.4]
  wire  _T_6726; // @[OneHot.scala 66:30:@3692.4]
  wire  _T_6727; // @[OneHot.scala 66:30:@3693.4]
  wire  _T_6728; // @[OneHot.scala 66:30:@3694.4]
  wire  _T_6729; // @[OneHot.scala 66:30:@3695.4]
  wire  _T_6730; // @[OneHot.scala 66:30:@3696.4]
  wire [15:0] _T_6771; // @[Mux.scala 31:69:@3714.4]
  wire [15:0] _T_6772; // @[Mux.scala 31:69:@3715.4]
  wire [15:0] _T_6773; // @[Mux.scala 31:69:@3716.4]
  wire [15:0] _T_6774; // @[Mux.scala 31:69:@3717.4]
  wire [15:0] _T_6775; // @[Mux.scala 31:69:@3718.4]
  wire [15:0] _T_6776; // @[Mux.scala 31:69:@3719.4]
  wire [15:0] _T_6777; // @[Mux.scala 31:69:@3720.4]
  wire [15:0] _T_6778; // @[Mux.scala 31:69:@3721.4]
  wire [15:0] _T_6779; // @[Mux.scala 31:69:@3722.4]
  wire [15:0] _T_6780; // @[Mux.scala 31:69:@3723.4]
  wire [15:0] _T_6781; // @[Mux.scala 31:69:@3724.4]
  wire [15:0] _T_6782; // @[Mux.scala 31:69:@3725.4]
  wire [15:0] _T_6783; // @[Mux.scala 31:69:@3726.4]
  wire [15:0] _T_6784; // @[Mux.scala 31:69:@3727.4]
  wire [15:0] _T_6785; // @[Mux.scala 31:69:@3728.4]
  wire [15:0] _T_6786; // @[Mux.scala 31:69:@3729.4]
  wire  _T_6787; // @[OneHot.scala 66:30:@3730.4]
  wire  _T_6788; // @[OneHot.scala 66:30:@3731.4]
  wire  _T_6789; // @[OneHot.scala 66:30:@3732.4]
  wire  _T_6790; // @[OneHot.scala 66:30:@3733.4]
  wire  _T_6791; // @[OneHot.scala 66:30:@3734.4]
  wire  _T_6792; // @[OneHot.scala 66:30:@3735.4]
  wire  _T_6793; // @[OneHot.scala 66:30:@3736.4]
  wire  _T_6794; // @[OneHot.scala 66:30:@3737.4]
  wire  _T_6795; // @[OneHot.scala 66:30:@3738.4]
  wire  _T_6796; // @[OneHot.scala 66:30:@3739.4]
  wire  _T_6797; // @[OneHot.scala 66:30:@3740.4]
  wire  _T_6798; // @[OneHot.scala 66:30:@3741.4]
  wire  _T_6799; // @[OneHot.scala 66:30:@3742.4]
  wire  _T_6800; // @[OneHot.scala 66:30:@3743.4]
  wire  _T_6801; // @[OneHot.scala 66:30:@3744.4]
  wire  _T_6802; // @[OneHot.scala 66:30:@3745.4]
  wire [15:0] _T_6843; // @[Mux.scala 31:69:@3763.4]
  wire [15:0] _T_6844; // @[Mux.scala 31:69:@3764.4]
  wire [15:0] _T_6845; // @[Mux.scala 31:69:@3765.4]
  wire [15:0] _T_6846; // @[Mux.scala 31:69:@3766.4]
  wire [15:0] _T_6847; // @[Mux.scala 31:69:@3767.4]
  wire [15:0] _T_6848; // @[Mux.scala 31:69:@3768.4]
  wire [15:0] _T_6849; // @[Mux.scala 31:69:@3769.4]
  wire [15:0] _T_6850; // @[Mux.scala 31:69:@3770.4]
  wire [15:0] _T_6851; // @[Mux.scala 31:69:@3771.4]
  wire [15:0] _T_6852; // @[Mux.scala 31:69:@3772.4]
  wire [15:0] _T_6853; // @[Mux.scala 31:69:@3773.4]
  wire [15:0] _T_6854; // @[Mux.scala 31:69:@3774.4]
  wire [15:0] _T_6855; // @[Mux.scala 31:69:@3775.4]
  wire [15:0] _T_6856; // @[Mux.scala 31:69:@3776.4]
  wire [15:0] _T_6857; // @[Mux.scala 31:69:@3777.4]
  wire [15:0] _T_6858; // @[Mux.scala 31:69:@3778.4]
  wire  _T_6859; // @[OneHot.scala 66:30:@3779.4]
  wire  _T_6860; // @[OneHot.scala 66:30:@3780.4]
  wire  _T_6861; // @[OneHot.scala 66:30:@3781.4]
  wire  _T_6862; // @[OneHot.scala 66:30:@3782.4]
  wire  _T_6863; // @[OneHot.scala 66:30:@3783.4]
  wire  _T_6864; // @[OneHot.scala 66:30:@3784.4]
  wire  _T_6865; // @[OneHot.scala 66:30:@3785.4]
  wire  _T_6866; // @[OneHot.scala 66:30:@3786.4]
  wire  _T_6867; // @[OneHot.scala 66:30:@3787.4]
  wire  _T_6868; // @[OneHot.scala 66:30:@3788.4]
  wire  _T_6869; // @[OneHot.scala 66:30:@3789.4]
  wire  _T_6870; // @[OneHot.scala 66:30:@3790.4]
  wire  _T_6871; // @[OneHot.scala 66:30:@3791.4]
  wire  _T_6872; // @[OneHot.scala 66:30:@3792.4]
  wire  _T_6873; // @[OneHot.scala 66:30:@3793.4]
  wire  _T_6874; // @[OneHot.scala 66:30:@3794.4]
  wire [15:0] _T_6915; // @[Mux.scala 31:69:@3812.4]
  wire [15:0] _T_6916; // @[Mux.scala 31:69:@3813.4]
  wire [15:0] _T_6917; // @[Mux.scala 31:69:@3814.4]
  wire [15:0] _T_6918; // @[Mux.scala 31:69:@3815.4]
  wire [15:0] _T_6919; // @[Mux.scala 31:69:@3816.4]
  wire [15:0] _T_6920; // @[Mux.scala 31:69:@3817.4]
  wire [15:0] _T_6921; // @[Mux.scala 31:69:@3818.4]
  wire [15:0] _T_6922; // @[Mux.scala 31:69:@3819.4]
  wire [15:0] _T_6923; // @[Mux.scala 31:69:@3820.4]
  wire [15:0] _T_6924; // @[Mux.scala 31:69:@3821.4]
  wire [15:0] _T_6925; // @[Mux.scala 31:69:@3822.4]
  wire [15:0] _T_6926; // @[Mux.scala 31:69:@3823.4]
  wire [15:0] _T_6927; // @[Mux.scala 31:69:@3824.4]
  wire [15:0] _T_6928; // @[Mux.scala 31:69:@3825.4]
  wire [15:0] _T_6929; // @[Mux.scala 31:69:@3826.4]
  wire [15:0] _T_6930; // @[Mux.scala 31:69:@3827.4]
  wire  _T_6931; // @[OneHot.scala 66:30:@3828.4]
  wire  _T_6932; // @[OneHot.scala 66:30:@3829.4]
  wire  _T_6933; // @[OneHot.scala 66:30:@3830.4]
  wire  _T_6934; // @[OneHot.scala 66:30:@3831.4]
  wire  _T_6935; // @[OneHot.scala 66:30:@3832.4]
  wire  _T_6936; // @[OneHot.scala 66:30:@3833.4]
  wire  _T_6937; // @[OneHot.scala 66:30:@3834.4]
  wire  _T_6938; // @[OneHot.scala 66:30:@3835.4]
  wire  _T_6939; // @[OneHot.scala 66:30:@3836.4]
  wire  _T_6940; // @[OneHot.scala 66:30:@3837.4]
  wire  _T_6941; // @[OneHot.scala 66:30:@3838.4]
  wire  _T_6942; // @[OneHot.scala 66:30:@3839.4]
  wire  _T_6943; // @[OneHot.scala 66:30:@3840.4]
  wire  _T_6944; // @[OneHot.scala 66:30:@3841.4]
  wire  _T_6945; // @[OneHot.scala 66:30:@3842.4]
  wire  _T_6946; // @[OneHot.scala 66:30:@3843.4]
  wire [15:0] _T_6987; // @[Mux.scala 31:69:@3861.4]
  wire [15:0] _T_6988; // @[Mux.scala 31:69:@3862.4]
  wire [15:0] _T_6989; // @[Mux.scala 31:69:@3863.4]
  wire [15:0] _T_6990; // @[Mux.scala 31:69:@3864.4]
  wire [15:0] _T_6991; // @[Mux.scala 31:69:@3865.4]
  wire [15:0] _T_6992; // @[Mux.scala 31:69:@3866.4]
  wire [15:0] _T_6993; // @[Mux.scala 31:69:@3867.4]
  wire [15:0] _T_6994; // @[Mux.scala 31:69:@3868.4]
  wire [15:0] _T_6995; // @[Mux.scala 31:69:@3869.4]
  wire [15:0] _T_6996; // @[Mux.scala 31:69:@3870.4]
  wire [15:0] _T_6997; // @[Mux.scala 31:69:@3871.4]
  wire [15:0] _T_6998; // @[Mux.scala 31:69:@3872.4]
  wire [15:0] _T_6999; // @[Mux.scala 31:69:@3873.4]
  wire [15:0] _T_7000; // @[Mux.scala 31:69:@3874.4]
  wire [15:0] _T_7001; // @[Mux.scala 31:69:@3875.4]
  wire [15:0] _T_7002; // @[Mux.scala 31:69:@3876.4]
  wire  _T_7003; // @[OneHot.scala 66:30:@3877.4]
  wire  _T_7004; // @[OneHot.scala 66:30:@3878.4]
  wire  _T_7005; // @[OneHot.scala 66:30:@3879.4]
  wire  _T_7006; // @[OneHot.scala 66:30:@3880.4]
  wire  _T_7007; // @[OneHot.scala 66:30:@3881.4]
  wire  _T_7008; // @[OneHot.scala 66:30:@3882.4]
  wire  _T_7009; // @[OneHot.scala 66:30:@3883.4]
  wire  _T_7010; // @[OneHot.scala 66:30:@3884.4]
  wire  _T_7011; // @[OneHot.scala 66:30:@3885.4]
  wire  _T_7012; // @[OneHot.scala 66:30:@3886.4]
  wire  _T_7013; // @[OneHot.scala 66:30:@3887.4]
  wire  _T_7014; // @[OneHot.scala 66:30:@3888.4]
  wire  _T_7015; // @[OneHot.scala 66:30:@3889.4]
  wire  _T_7016; // @[OneHot.scala 66:30:@3890.4]
  wire  _T_7017; // @[OneHot.scala 66:30:@3891.4]
  wire  _T_7018; // @[OneHot.scala 66:30:@3892.4]
  wire [15:0] _T_7059; // @[Mux.scala 31:69:@3910.4]
  wire [15:0] _T_7060; // @[Mux.scala 31:69:@3911.4]
  wire [15:0] _T_7061; // @[Mux.scala 31:69:@3912.4]
  wire [15:0] _T_7062; // @[Mux.scala 31:69:@3913.4]
  wire [15:0] _T_7063; // @[Mux.scala 31:69:@3914.4]
  wire [15:0] _T_7064; // @[Mux.scala 31:69:@3915.4]
  wire [15:0] _T_7065; // @[Mux.scala 31:69:@3916.4]
  wire [15:0] _T_7066; // @[Mux.scala 31:69:@3917.4]
  wire [15:0] _T_7067; // @[Mux.scala 31:69:@3918.4]
  wire [15:0] _T_7068; // @[Mux.scala 31:69:@3919.4]
  wire [15:0] _T_7069; // @[Mux.scala 31:69:@3920.4]
  wire [15:0] _T_7070; // @[Mux.scala 31:69:@3921.4]
  wire [15:0] _T_7071; // @[Mux.scala 31:69:@3922.4]
  wire [15:0] _T_7072; // @[Mux.scala 31:69:@3923.4]
  wire [15:0] _T_7073; // @[Mux.scala 31:69:@3924.4]
  wire [15:0] _T_7074; // @[Mux.scala 31:69:@3925.4]
  wire  _T_7075; // @[OneHot.scala 66:30:@3926.4]
  wire  _T_7076; // @[OneHot.scala 66:30:@3927.4]
  wire  _T_7077; // @[OneHot.scala 66:30:@3928.4]
  wire  _T_7078; // @[OneHot.scala 66:30:@3929.4]
  wire  _T_7079; // @[OneHot.scala 66:30:@3930.4]
  wire  _T_7080; // @[OneHot.scala 66:30:@3931.4]
  wire  _T_7081; // @[OneHot.scala 66:30:@3932.4]
  wire  _T_7082; // @[OneHot.scala 66:30:@3933.4]
  wire  _T_7083; // @[OneHot.scala 66:30:@3934.4]
  wire  _T_7084; // @[OneHot.scala 66:30:@3935.4]
  wire  _T_7085; // @[OneHot.scala 66:30:@3936.4]
  wire  _T_7086; // @[OneHot.scala 66:30:@3937.4]
  wire  _T_7087; // @[OneHot.scala 66:30:@3938.4]
  wire  _T_7088; // @[OneHot.scala 66:30:@3939.4]
  wire  _T_7089; // @[OneHot.scala 66:30:@3940.4]
  wire  _T_7090; // @[OneHot.scala 66:30:@3941.4]
  wire [7:0] _T_7155; // @[Mux.scala 19:72:@3965.4]
  wire [15:0] _T_7163; // @[Mux.scala 19:72:@3973.4]
  wire [15:0] _T_7165; // @[Mux.scala 19:72:@3974.4]
  wire [7:0] _T_7172; // @[Mux.scala 19:72:@3981.4]
  wire [15:0] _T_7180; // @[Mux.scala 19:72:@3989.4]
  wire [15:0] _T_7182; // @[Mux.scala 19:72:@3990.4]
  wire [7:0] _T_7189; // @[Mux.scala 19:72:@3997.4]
  wire [15:0] _T_7197; // @[Mux.scala 19:72:@4005.4]
  wire [15:0] _T_7199; // @[Mux.scala 19:72:@4006.4]
  wire [7:0] _T_7206; // @[Mux.scala 19:72:@4013.4]
  wire [15:0] _T_7214; // @[Mux.scala 19:72:@4021.4]
  wire [15:0] _T_7216; // @[Mux.scala 19:72:@4022.4]
  wire [7:0] _T_7223; // @[Mux.scala 19:72:@4029.4]
  wire [15:0] _T_7231; // @[Mux.scala 19:72:@4037.4]
  wire [15:0] _T_7233; // @[Mux.scala 19:72:@4038.4]
  wire [7:0] _T_7240; // @[Mux.scala 19:72:@4045.4]
  wire [15:0] _T_7248; // @[Mux.scala 19:72:@4053.4]
  wire [15:0] _T_7250; // @[Mux.scala 19:72:@4054.4]
  wire [7:0] _T_7257; // @[Mux.scala 19:72:@4061.4]
  wire [15:0] _T_7265; // @[Mux.scala 19:72:@4069.4]
  wire [15:0] _T_7267; // @[Mux.scala 19:72:@4070.4]
  wire [7:0] _T_7274; // @[Mux.scala 19:72:@4077.4]
  wire [15:0] _T_7282; // @[Mux.scala 19:72:@4085.4]
  wire [15:0] _T_7284; // @[Mux.scala 19:72:@4086.4]
  wire [7:0] _T_7291; // @[Mux.scala 19:72:@4093.4]
  wire [15:0] _T_7299; // @[Mux.scala 19:72:@4101.4]
  wire [15:0] _T_7301; // @[Mux.scala 19:72:@4102.4]
  wire [7:0] _T_7308; // @[Mux.scala 19:72:@4109.4]
  wire [15:0] _T_7316; // @[Mux.scala 19:72:@4117.4]
  wire [15:0] _T_7318; // @[Mux.scala 19:72:@4118.4]
  wire [7:0] _T_7325; // @[Mux.scala 19:72:@4125.4]
  wire [15:0] _T_7333; // @[Mux.scala 19:72:@4133.4]
  wire [15:0] _T_7335; // @[Mux.scala 19:72:@4134.4]
  wire [7:0] _T_7342; // @[Mux.scala 19:72:@4141.4]
  wire [15:0] _T_7350; // @[Mux.scala 19:72:@4149.4]
  wire [15:0] _T_7352; // @[Mux.scala 19:72:@4150.4]
  wire [7:0] _T_7359; // @[Mux.scala 19:72:@4157.4]
  wire [15:0] _T_7367; // @[Mux.scala 19:72:@4165.4]
  wire [15:0] _T_7369; // @[Mux.scala 19:72:@4166.4]
  wire [7:0] _T_7376; // @[Mux.scala 19:72:@4173.4]
  wire [15:0] _T_7384; // @[Mux.scala 19:72:@4181.4]
  wire [15:0] _T_7386; // @[Mux.scala 19:72:@4182.4]
  wire [7:0] _T_7393; // @[Mux.scala 19:72:@4189.4]
  wire [15:0] _T_7401; // @[Mux.scala 19:72:@4197.4]
  wire [15:0] _T_7403; // @[Mux.scala 19:72:@4198.4]
  wire [7:0] _T_7410; // @[Mux.scala 19:72:@4205.4]
  wire [15:0] _T_7418; // @[Mux.scala 19:72:@4213.4]
  wire [15:0] _T_7420; // @[Mux.scala 19:72:@4214.4]
  wire [15:0] _T_7421; // @[Mux.scala 19:72:@4215.4]
  wire [15:0] _T_7422; // @[Mux.scala 19:72:@4216.4]
  wire [15:0] _T_7423; // @[Mux.scala 19:72:@4217.4]
  wire [15:0] _T_7424; // @[Mux.scala 19:72:@4218.4]
  wire [15:0] _T_7425; // @[Mux.scala 19:72:@4219.4]
  wire [15:0] _T_7426; // @[Mux.scala 19:72:@4220.4]
  wire [15:0] _T_7427; // @[Mux.scala 19:72:@4221.4]
  wire [15:0] _T_7428; // @[Mux.scala 19:72:@4222.4]
  wire [15:0] _T_7429; // @[Mux.scala 19:72:@4223.4]
  wire [15:0] _T_7430; // @[Mux.scala 19:72:@4224.4]
  wire [15:0] _T_7431; // @[Mux.scala 19:72:@4225.4]
  wire [15:0] _T_7432; // @[Mux.scala 19:72:@4226.4]
  wire [15:0] _T_7433; // @[Mux.scala 19:72:@4227.4]
  wire [15:0] _T_7434; // @[Mux.scala 19:72:@4228.4]
  wire [15:0] _T_7435; // @[Mux.scala 19:72:@4229.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@4233.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@4235.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@4237.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@4239.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@4241.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@4243.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@4245.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@4247.4]
  wire  inputDataPriorityPorts_0_8; // @[Mux.scala 19:72:@4249.4]
  wire  inputDataPriorityPorts_0_9; // @[Mux.scala 19:72:@4251.4]
  wire  inputDataPriorityPorts_0_10; // @[Mux.scala 19:72:@4253.4]
  wire  inputDataPriorityPorts_0_11; // @[Mux.scala 19:72:@4255.4]
  wire  inputDataPriorityPorts_0_12; // @[Mux.scala 19:72:@4257.4]
  wire  inputDataPriorityPorts_0_13; // @[Mux.scala 19:72:@4259.4]
  wire  inputDataPriorityPorts_0_14; // @[Mux.scala 19:72:@4261.4]
  wire  inputDataPriorityPorts_0_15; // @[Mux.scala 19:72:@4263.4]
  wire  _T_7581; // @[StoreQueue.scala 209:52:@4287.6]
  wire  _T_7582; // @[StoreQueue.scala 209:81:@4288.6]
  wire [31:0] _GEN_992; // @[StoreQueue.scala 210:40:@4292.6]
  wire  _GEN_993; // @[StoreQueue.scala 210:40:@4292.6]
  wire  _T_7598; // @[StoreQueue.scala 215:52:@4297.6]
  wire  _T_7599; // @[StoreQueue.scala 215:81:@4298.6]
  wire [31:0] _GEN_994; // @[StoreQueue.scala 216:40:@4302.6]
  wire  _GEN_995; // @[StoreQueue.scala 216:40:@4302.6]
  wire  _GEN_996; // @[StoreQueue.scala 204:35:@4281.4]
  wire  _GEN_997; // @[StoreQueue.scala 204:35:@4281.4]
  wire [31:0] _GEN_998; // @[StoreQueue.scala 204:35:@4281.4]
  wire [31:0] _GEN_999; // @[StoreQueue.scala 204:35:@4281.4]
  wire  _T_7617; // @[StoreQueue.scala 209:52:@4313.6]
  wire  _T_7618; // @[StoreQueue.scala 209:81:@4314.6]
  wire [31:0] _GEN_1000; // @[StoreQueue.scala 210:40:@4318.6]
  wire  _GEN_1001; // @[StoreQueue.scala 210:40:@4318.6]
  wire  _T_7634; // @[StoreQueue.scala 215:52:@4323.6]
  wire  _T_7635; // @[StoreQueue.scala 215:81:@4324.6]
  wire [31:0] _GEN_1002; // @[StoreQueue.scala 216:40:@4328.6]
  wire  _GEN_1003; // @[StoreQueue.scala 216:40:@4328.6]
  wire  _GEN_1004; // @[StoreQueue.scala 204:35:@4307.4]
  wire  _GEN_1005; // @[StoreQueue.scala 204:35:@4307.4]
  wire [31:0] _GEN_1006; // @[StoreQueue.scala 204:35:@4307.4]
  wire [31:0] _GEN_1007; // @[StoreQueue.scala 204:35:@4307.4]
  wire  _T_7653; // @[StoreQueue.scala 209:52:@4339.6]
  wire  _T_7654; // @[StoreQueue.scala 209:81:@4340.6]
  wire [31:0] _GEN_1008; // @[StoreQueue.scala 210:40:@4344.6]
  wire  _GEN_1009; // @[StoreQueue.scala 210:40:@4344.6]
  wire  _T_7670; // @[StoreQueue.scala 215:52:@4349.6]
  wire  _T_7671; // @[StoreQueue.scala 215:81:@4350.6]
  wire [31:0] _GEN_1010; // @[StoreQueue.scala 216:40:@4354.6]
  wire  _GEN_1011; // @[StoreQueue.scala 216:40:@4354.6]
  wire  _GEN_1012; // @[StoreQueue.scala 204:35:@4333.4]
  wire  _GEN_1013; // @[StoreQueue.scala 204:35:@4333.4]
  wire [31:0] _GEN_1014; // @[StoreQueue.scala 204:35:@4333.4]
  wire [31:0] _GEN_1015; // @[StoreQueue.scala 204:35:@4333.4]
  wire  _T_7689; // @[StoreQueue.scala 209:52:@4365.6]
  wire  _T_7690; // @[StoreQueue.scala 209:81:@4366.6]
  wire [31:0] _GEN_1016; // @[StoreQueue.scala 210:40:@4370.6]
  wire  _GEN_1017; // @[StoreQueue.scala 210:40:@4370.6]
  wire  _T_7706; // @[StoreQueue.scala 215:52:@4375.6]
  wire  _T_7707; // @[StoreQueue.scala 215:81:@4376.6]
  wire [31:0] _GEN_1018; // @[StoreQueue.scala 216:40:@4380.6]
  wire  _GEN_1019; // @[StoreQueue.scala 216:40:@4380.6]
  wire  _GEN_1020; // @[StoreQueue.scala 204:35:@4359.4]
  wire  _GEN_1021; // @[StoreQueue.scala 204:35:@4359.4]
  wire [31:0] _GEN_1022; // @[StoreQueue.scala 204:35:@4359.4]
  wire [31:0] _GEN_1023; // @[StoreQueue.scala 204:35:@4359.4]
  wire  _T_7725; // @[StoreQueue.scala 209:52:@4391.6]
  wire  _T_7726; // @[StoreQueue.scala 209:81:@4392.6]
  wire [31:0] _GEN_1024; // @[StoreQueue.scala 210:40:@4396.6]
  wire  _GEN_1025; // @[StoreQueue.scala 210:40:@4396.6]
  wire  _T_7742; // @[StoreQueue.scala 215:52:@4401.6]
  wire  _T_7743; // @[StoreQueue.scala 215:81:@4402.6]
  wire [31:0] _GEN_1026; // @[StoreQueue.scala 216:40:@4406.6]
  wire  _GEN_1027; // @[StoreQueue.scala 216:40:@4406.6]
  wire  _GEN_1028; // @[StoreQueue.scala 204:35:@4385.4]
  wire  _GEN_1029; // @[StoreQueue.scala 204:35:@4385.4]
  wire [31:0] _GEN_1030; // @[StoreQueue.scala 204:35:@4385.4]
  wire [31:0] _GEN_1031; // @[StoreQueue.scala 204:35:@4385.4]
  wire  _T_7761; // @[StoreQueue.scala 209:52:@4417.6]
  wire  _T_7762; // @[StoreQueue.scala 209:81:@4418.6]
  wire [31:0] _GEN_1032; // @[StoreQueue.scala 210:40:@4422.6]
  wire  _GEN_1033; // @[StoreQueue.scala 210:40:@4422.6]
  wire  _T_7778; // @[StoreQueue.scala 215:52:@4427.6]
  wire  _T_7779; // @[StoreQueue.scala 215:81:@4428.6]
  wire [31:0] _GEN_1034; // @[StoreQueue.scala 216:40:@4432.6]
  wire  _GEN_1035; // @[StoreQueue.scala 216:40:@4432.6]
  wire  _GEN_1036; // @[StoreQueue.scala 204:35:@4411.4]
  wire  _GEN_1037; // @[StoreQueue.scala 204:35:@4411.4]
  wire [31:0] _GEN_1038; // @[StoreQueue.scala 204:35:@4411.4]
  wire [31:0] _GEN_1039; // @[StoreQueue.scala 204:35:@4411.4]
  wire  _T_7797; // @[StoreQueue.scala 209:52:@4443.6]
  wire  _T_7798; // @[StoreQueue.scala 209:81:@4444.6]
  wire [31:0] _GEN_1040; // @[StoreQueue.scala 210:40:@4448.6]
  wire  _GEN_1041; // @[StoreQueue.scala 210:40:@4448.6]
  wire  _T_7814; // @[StoreQueue.scala 215:52:@4453.6]
  wire  _T_7815; // @[StoreQueue.scala 215:81:@4454.6]
  wire [31:0] _GEN_1042; // @[StoreQueue.scala 216:40:@4458.6]
  wire  _GEN_1043; // @[StoreQueue.scala 216:40:@4458.6]
  wire  _GEN_1044; // @[StoreQueue.scala 204:35:@4437.4]
  wire  _GEN_1045; // @[StoreQueue.scala 204:35:@4437.4]
  wire [31:0] _GEN_1046; // @[StoreQueue.scala 204:35:@4437.4]
  wire [31:0] _GEN_1047; // @[StoreQueue.scala 204:35:@4437.4]
  wire  _T_7833; // @[StoreQueue.scala 209:52:@4469.6]
  wire  _T_7834; // @[StoreQueue.scala 209:81:@4470.6]
  wire [31:0] _GEN_1048; // @[StoreQueue.scala 210:40:@4474.6]
  wire  _GEN_1049; // @[StoreQueue.scala 210:40:@4474.6]
  wire  _T_7850; // @[StoreQueue.scala 215:52:@4479.6]
  wire  _T_7851; // @[StoreQueue.scala 215:81:@4480.6]
  wire [31:0] _GEN_1050; // @[StoreQueue.scala 216:40:@4484.6]
  wire  _GEN_1051; // @[StoreQueue.scala 216:40:@4484.6]
  wire  _GEN_1052; // @[StoreQueue.scala 204:35:@4463.4]
  wire  _GEN_1053; // @[StoreQueue.scala 204:35:@4463.4]
  wire [31:0] _GEN_1054; // @[StoreQueue.scala 204:35:@4463.4]
  wire [31:0] _GEN_1055; // @[StoreQueue.scala 204:35:@4463.4]
  wire  _T_7869; // @[StoreQueue.scala 209:52:@4495.6]
  wire  _T_7870; // @[StoreQueue.scala 209:81:@4496.6]
  wire [31:0] _GEN_1056; // @[StoreQueue.scala 210:40:@4500.6]
  wire  _GEN_1057; // @[StoreQueue.scala 210:40:@4500.6]
  wire  _T_7886; // @[StoreQueue.scala 215:52:@4505.6]
  wire  _T_7887; // @[StoreQueue.scala 215:81:@4506.6]
  wire [31:0] _GEN_1058; // @[StoreQueue.scala 216:40:@4510.6]
  wire  _GEN_1059; // @[StoreQueue.scala 216:40:@4510.6]
  wire  _GEN_1060; // @[StoreQueue.scala 204:35:@4489.4]
  wire  _GEN_1061; // @[StoreQueue.scala 204:35:@4489.4]
  wire [31:0] _GEN_1062; // @[StoreQueue.scala 204:35:@4489.4]
  wire [31:0] _GEN_1063; // @[StoreQueue.scala 204:35:@4489.4]
  wire  _T_7905; // @[StoreQueue.scala 209:52:@4521.6]
  wire  _T_7906; // @[StoreQueue.scala 209:81:@4522.6]
  wire [31:0] _GEN_1064; // @[StoreQueue.scala 210:40:@4526.6]
  wire  _GEN_1065; // @[StoreQueue.scala 210:40:@4526.6]
  wire  _T_7922; // @[StoreQueue.scala 215:52:@4531.6]
  wire  _T_7923; // @[StoreQueue.scala 215:81:@4532.6]
  wire [31:0] _GEN_1066; // @[StoreQueue.scala 216:40:@4536.6]
  wire  _GEN_1067; // @[StoreQueue.scala 216:40:@4536.6]
  wire  _GEN_1068; // @[StoreQueue.scala 204:35:@4515.4]
  wire  _GEN_1069; // @[StoreQueue.scala 204:35:@4515.4]
  wire [31:0] _GEN_1070; // @[StoreQueue.scala 204:35:@4515.4]
  wire [31:0] _GEN_1071; // @[StoreQueue.scala 204:35:@4515.4]
  wire  _T_7941; // @[StoreQueue.scala 209:52:@4547.6]
  wire  _T_7942; // @[StoreQueue.scala 209:81:@4548.6]
  wire [31:0] _GEN_1072; // @[StoreQueue.scala 210:40:@4552.6]
  wire  _GEN_1073; // @[StoreQueue.scala 210:40:@4552.6]
  wire  _T_7958; // @[StoreQueue.scala 215:52:@4557.6]
  wire  _T_7959; // @[StoreQueue.scala 215:81:@4558.6]
  wire [31:0] _GEN_1074; // @[StoreQueue.scala 216:40:@4562.6]
  wire  _GEN_1075; // @[StoreQueue.scala 216:40:@4562.6]
  wire  _GEN_1076; // @[StoreQueue.scala 204:35:@4541.4]
  wire  _GEN_1077; // @[StoreQueue.scala 204:35:@4541.4]
  wire [31:0] _GEN_1078; // @[StoreQueue.scala 204:35:@4541.4]
  wire [31:0] _GEN_1079; // @[StoreQueue.scala 204:35:@4541.4]
  wire  _T_7977; // @[StoreQueue.scala 209:52:@4573.6]
  wire  _T_7978; // @[StoreQueue.scala 209:81:@4574.6]
  wire [31:0] _GEN_1080; // @[StoreQueue.scala 210:40:@4578.6]
  wire  _GEN_1081; // @[StoreQueue.scala 210:40:@4578.6]
  wire  _T_7994; // @[StoreQueue.scala 215:52:@4583.6]
  wire  _T_7995; // @[StoreQueue.scala 215:81:@4584.6]
  wire [31:0] _GEN_1082; // @[StoreQueue.scala 216:40:@4588.6]
  wire  _GEN_1083; // @[StoreQueue.scala 216:40:@4588.6]
  wire  _GEN_1084; // @[StoreQueue.scala 204:35:@4567.4]
  wire  _GEN_1085; // @[StoreQueue.scala 204:35:@4567.4]
  wire [31:0] _GEN_1086; // @[StoreQueue.scala 204:35:@4567.4]
  wire [31:0] _GEN_1087; // @[StoreQueue.scala 204:35:@4567.4]
  wire  _T_8013; // @[StoreQueue.scala 209:52:@4599.6]
  wire  _T_8014; // @[StoreQueue.scala 209:81:@4600.6]
  wire [31:0] _GEN_1088; // @[StoreQueue.scala 210:40:@4604.6]
  wire  _GEN_1089; // @[StoreQueue.scala 210:40:@4604.6]
  wire  _T_8030; // @[StoreQueue.scala 215:52:@4609.6]
  wire  _T_8031; // @[StoreQueue.scala 215:81:@4610.6]
  wire [31:0] _GEN_1090; // @[StoreQueue.scala 216:40:@4614.6]
  wire  _GEN_1091; // @[StoreQueue.scala 216:40:@4614.6]
  wire  _GEN_1092; // @[StoreQueue.scala 204:35:@4593.4]
  wire  _GEN_1093; // @[StoreQueue.scala 204:35:@4593.4]
  wire [31:0] _GEN_1094; // @[StoreQueue.scala 204:35:@4593.4]
  wire [31:0] _GEN_1095; // @[StoreQueue.scala 204:35:@4593.4]
  wire  _T_8049; // @[StoreQueue.scala 209:52:@4625.6]
  wire  _T_8050; // @[StoreQueue.scala 209:81:@4626.6]
  wire [31:0] _GEN_1096; // @[StoreQueue.scala 210:40:@4630.6]
  wire  _GEN_1097; // @[StoreQueue.scala 210:40:@4630.6]
  wire  _T_8066; // @[StoreQueue.scala 215:52:@4635.6]
  wire  _T_8067; // @[StoreQueue.scala 215:81:@4636.6]
  wire [31:0] _GEN_1098; // @[StoreQueue.scala 216:40:@4640.6]
  wire  _GEN_1099; // @[StoreQueue.scala 216:40:@4640.6]
  wire  _GEN_1100; // @[StoreQueue.scala 204:35:@4619.4]
  wire  _GEN_1101; // @[StoreQueue.scala 204:35:@4619.4]
  wire [31:0] _GEN_1102; // @[StoreQueue.scala 204:35:@4619.4]
  wire [31:0] _GEN_1103; // @[StoreQueue.scala 204:35:@4619.4]
  wire  _T_8085; // @[StoreQueue.scala 209:52:@4651.6]
  wire  _T_8086; // @[StoreQueue.scala 209:81:@4652.6]
  wire [31:0] _GEN_1104; // @[StoreQueue.scala 210:40:@4656.6]
  wire  _GEN_1105; // @[StoreQueue.scala 210:40:@4656.6]
  wire  _T_8102; // @[StoreQueue.scala 215:52:@4661.6]
  wire  _T_8103; // @[StoreQueue.scala 215:81:@4662.6]
  wire [31:0] _GEN_1106; // @[StoreQueue.scala 216:40:@4666.6]
  wire  _GEN_1107; // @[StoreQueue.scala 216:40:@4666.6]
  wire  _GEN_1108; // @[StoreQueue.scala 204:35:@4645.4]
  wire  _GEN_1109; // @[StoreQueue.scala 204:35:@4645.4]
  wire [31:0] _GEN_1110; // @[StoreQueue.scala 204:35:@4645.4]
  wire [31:0] _GEN_1111; // @[StoreQueue.scala 204:35:@4645.4]
  wire  _T_8121; // @[StoreQueue.scala 209:52:@4677.6]
  wire  _T_8122; // @[StoreQueue.scala 209:81:@4678.6]
  wire [31:0] _GEN_1112; // @[StoreQueue.scala 210:40:@4682.6]
  wire  _GEN_1113; // @[StoreQueue.scala 210:40:@4682.6]
  wire  _T_8138; // @[StoreQueue.scala 215:52:@4687.6]
  wire  _T_8139; // @[StoreQueue.scala 215:81:@4688.6]
  wire [31:0] _GEN_1114; // @[StoreQueue.scala 216:40:@4692.6]
  wire  _GEN_1115; // @[StoreQueue.scala 216:40:@4692.6]
  wire  _GEN_1116; // @[StoreQueue.scala 204:35:@4671.4]
  wire  _GEN_1117; // @[StoreQueue.scala 204:35:@4671.4]
  wire [31:0] _GEN_1118; // @[StoreQueue.scala 204:35:@4671.4]
  wire [31:0] _GEN_1119; // @[StoreQueue.scala 204:35:@4671.4]
  wire  _T_8153; // @[StoreQueue.scala 229:23:@4697.4]
  wire [4:0] _T_8156; // @[util.scala 10:8:@4699.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@4700.6]
  wire [4:0] _T_8157; // @[util.scala 10:14:@4700.6]
  wire [4:0] _GEN_1120; // @[StoreQueue.scala 229:50:@4698.4]
  wire [3:0] _GEN_1234; // @[util.scala 10:8:@4704.6]
  wire [4:0] _T_8159; // @[util.scala 10:8:@4704.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@4705.6]
  wire [4:0] _T_8160; // @[util.scala 10:14:@4705.6]
  wire [4:0] _GEN_1121; // @[StoreQueue.scala 233:20:@4703.4]
  wire  _T_8162; // @[StoreQueue.scala 237:84:@4708.4]
  wire  _T_8163; // @[StoreQueue.scala 237:81:@4709.4]
  wire  _T_8165; // @[StoreQueue.scala 237:84:@4710.4]
  wire  _T_8166; // @[StoreQueue.scala 237:81:@4711.4]
  wire  _T_8168; // @[StoreQueue.scala 237:84:@4712.4]
  wire  _T_8169; // @[StoreQueue.scala 237:81:@4713.4]
  wire  _T_8171; // @[StoreQueue.scala 237:84:@4714.4]
  wire  _T_8172; // @[StoreQueue.scala 237:81:@4715.4]
  wire  _T_8174; // @[StoreQueue.scala 237:84:@4716.4]
  wire  _T_8175; // @[StoreQueue.scala 237:81:@4717.4]
  wire  _T_8177; // @[StoreQueue.scala 237:84:@4718.4]
  wire  _T_8178; // @[StoreQueue.scala 237:81:@4719.4]
  wire  _T_8180; // @[StoreQueue.scala 237:84:@4720.4]
  wire  _T_8181; // @[StoreQueue.scala 237:81:@4721.4]
  wire  _T_8183; // @[StoreQueue.scala 237:84:@4722.4]
  wire  _T_8184; // @[StoreQueue.scala 237:81:@4723.4]
  wire  _T_8186; // @[StoreQueue.scala 237:84:@4724.4]
  wire  _T_8187; // @[StoreQueue.scala 237:81:@4725.4]
  wire  _T_8189; // @[StoreQueue.scala 237:84:@4726.4]
  wire  _T_8190; // @[StoreQueue.scala 237:81:@4727.4]
  wire  _T_8192; // @[StoreQueue.scala 237:84:@4728.4]
  wire  _T_8193; // @[StoreQueue.scala 237:81:@4729.4]
  wire  _T_8195; // @[StoreQueue.scala 237:84:@4730.4]
  wire  _T_8196; // @[StoreQueue.scala 237:81:@4731.4]
  wire  _T_8198; // @[StoreQueue.scala 237:84:@4732.4]
  wire  _T_8199; // @[StoreQueue.scala 237:81:@4733.4]
  wire  _T_8201; // @[StoreQueue.scala 237:84:@4734.4]
  wire  _T_8202; // @[StoreQueue.scala 237:81:@4735.4]
  wire  _T_8204; // @[StoreQueue.scala 237:84:@4736.4]
  wire  _T_8205; // @[StoreQueue.scala 237:81:@4737.4]
  wire  _T_8207; // @[StoreQueue.scala 237:84:@4738.4]
  wire  _T_8208; // @[StoreQueue.scala 237:81:@4739.4]
  wire  _T_8233; // @[StoreQueue.scala 237:98:@4758.4]
  wire  _T_8234; // @[StoreQueue.scala 237:98:@4759.4]
  wire  _T_8235; // @[StoreQueue.scala 237:98:@4760.4]
  wire  _T_8236; // @[StoreQueue.scala 237:98:@4761.4]
  wire  _T_8237; // @[StoreQueue.scala 237:98:@4762.4]
  wire  _T_8238; // @[StoreQueue.scala 237:98:@4763.4]
  wire  _T_8239; // @[StoreQueue.scala 237:98:@4764.4]
  wire  _T_8240; // @[StoreQueue.scala 237:98:@4765.4]
  wire  _T_8241; // @[StoreQueue.scala 237:98:@4766.4]
  wire  _T_8242; // @[StoreQueue.scala 237:98:@4767.4]
  wire  _T_8243; // @[StoreQueue.scala 237:98:@4768.4]
  wire  _T_8244; // @[StoreQueue.scala 237:98:@4769.4]
  wire  _T_8245; // @[StoreQueue.scala 237:98:@4770.4]
  wire  _T_8246; // @[StoreQueue.scala 237:98:@4771.4]
  wire [31:0] _GEN_1123; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1124; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1125; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1126; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1127; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1128; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1129; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1130; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1131; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1132; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1133; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1134; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1135; // @[StoreQueue.scala 252:21:@4841.4]
  wire [31:0] _GEN_1136; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1138 = {{2'd0}, tail}; // @[util.scala 14:20:@173.4]
  assign _T_1596 = 6'h10 - _GEN_1138; // @[util.scala 14:20:@173.4]
  assign _T_1597 = $unsigned(_T_1596); // @[util.scala 14:20:@174.4]
  assign _T_1598 = _T_1597[5:0]; // @[util.scala 14:20:@175.4]
  assign _GEN_0 = _T_1598 % 6'h10; // @[util.scala 14:25:@176.4]
  assign _T_1599 = _GEN_0[4:0]; // @[util.scala 14:25:@176.4]
  assign _GEN_1139 = {{4'd0}, io_bbNumStores}; // @[StoreQueue.scala 70:46:@177.4]
  assign _T_1600 = _T_1599 < _GEN_1139; // @[StoreQueue.scala 70:46:@177.4]
  assign initBits_0 = _T_1600 & io_bbStart; // @[StoreQueue.scala 70:64:@178.4]
  assign _T_1605 = 6'h11 - _GEN_1138; // @[util.scala 14:20:@180.4]
  assign _T_1606 = $unsigned(_T_1605); // @[util.scala 14:20:@181.4]
  assign _T_1607 = _T_1606[5:0]; // @[util.scala 14:20:@182.4]
  assign _GEN_16 = _T_1607 % 6'h10; // @[util.scala 14:25:@183.4]
  assign _T_1608 = _GEN_16[4:0]; // @[util.scala 14:25:@183.4]
  assign _T_1609 = _T_1608 < _GEN_1139; // @[StoreQueue.scala 70:46:@184.4]
  assign initBits_1 = _T_1609 & io_bbStart; // @[StoreQueue.scala 70:64:@185.4]
  assign _T_1614 = 6'h12 - _GEN_1138; // @[util.scala 14:20:@187.4]
  assign _T_1615 = $unsigned(_T_1614); // @[util.scala 14:20:@188.4]
  assign _T_1616 = _T_1615[5:0]; // @[util.scala 14:20:@189.4]
  assign _GEN_17 = _T_1616 % 6'h10; // @[util.scala 14:25:@190.4]
  assign _T_1617 = _GEN_17[4:0]; // @[util.scala 14:25:@190.4]
  assign _T_1618 = _T_1617 < _GEN_1139; // @[StoreQueue.scala 70:46:@191.4]
  assign initBits_2 = _T_1618 & io_bbStart; // @[StoreQueue.scala 70:64:@192.4]
  assign _T_1623 = 6'h13 - _GEN_1138; // @[util.scala 14:20:@194.4]
  assign _T_1624 = $unsigned(_T_1623); // @[util.scala 14:20:@195.4]
  assign _T_1625 = _T_1624[5:0]; // @[util.scala 14:20:@196.4]
  assign _GEN_18 = _T_1625 % 6'h10; // @[util.scala 14:25:@197.4]
  assign _T_1626 = _GEN_18[4:0]; // @[util.scala 14:25:@197.4]
  assign _T_1627 = _T_1626 < _GEN_1139; // @[StoreQueue.scala 70:46:@198.4]
  assign initBits_3 = _T_1627 & io_bbStart; // @[StoreQueue.scala 70:64:@199.4]
  assign _T_1632 = 6'h14 - _GEN_1138; // @[util.scala 14:20:@201.4]
  assign _T_1633 = $unsigned(_T_1632); // @[util.scala 14:20:@202.4]
  assign _T_1634 = _T_1633[5:0]; // @[util.scala 14:20:@203.4]
  assign _GEN_19 = _T_1634 % 6'h10; // @[util.scala 14:25:@204.4]
  assign _T_1635 = _GEN_19[4:0]; // @[util.scala 14:25:@204.4]
  assign _T_1636 = _T_1635 < _GEN_1139; // @[StoreQueue.scala 70:46:@205.4]
  assign initBits_4 = _T_1636 & io_bbStart; // @[StoreQueue.scala 70:64:@206.4]
  assign _T_1641 = 6'h15 - _GEN_1138; // @[util.scala 14:20:@208.4]
  assign _T_1642 = $unsigned(_T_1641); // @[util.scala 14:20:@209.4]
  assign _T_1643 = _T_1642[5:0]; // @[util.scala 14:20:@210.4]
  assign _GEN_20 = _T_1643 % 6'h10; // @[util.scala 14:25:@211.4]
  assign _T_1644 = _GEN_20[4:0]; // @[util.scala 14:25:@211.4]
  assign _T_1645 = _T_1644 < _GEN_1139; // @[StoreQueue.scala 70:46:@212.4]
  assign initBits_5 = _T_1645 & io_bbStart; // @[StoreQueue.scala 70:64:@213.4]
  assign _T_1650 = 6'h16 - _GEN_1138; // @[util.scala 14:20:@215.4]
  assign _T_1651 = $unsigned(_T_1650); // @[util.scala 14:20:@216.4]
  assign _T_1652 = _T_1651[5:0]; // @[util.scala 14:20:@217.4]
  assign _GEN_21 = _T_1652 % 6'h10; // @[util.scala 14:25:@218.4]
  assign _T_1653 = _GEN_21[4:0]; // @[util.scala 14:25:@218.4]
  assign _T_1654 = _T_1653 < _GEN_1139; // @[StoreQueue.scala 70:46:@219.4]
  assign initBits_6 = _T_1654 & io_bbStart; // @[StoreQueue.scala 70:64:@220.4]
  assign _T_1659 = 6'h17 - _GEN_1138; // @[util.scala 14:20:@222.4]
  assign _T_1660 = $unsigned(_T_1659); // @[util.scala 14:20:@223.4]
  assign _T_1661 = _T_1660[5:0]; // @[util.scala 14:20:@224.4]
  assign _GEN_22 = _T_1661 % 6'h10; // @[util.scala 14:25:@225.4]
  assign _T_1662 = _GEN_22[4:0]; // @[util.scala 14:25:@225.4]
  assign _T_1663 = _T_1662 < _GEN_1139; // @[StoreQueue.scala 70:46:@226.4]
  assign initBits_7 = _T_1663 & io_bbStart; // @[StoreQueue.scala 70:64:@227.4]
  assign _T_1668 = 6'h18 - _GEN_1138; // @[util.scala 14:20:@229.4]
  assign _T_1669 = $unsigned(_T_1668); // @[util.scala 14:20:@230.4]
  assign _T_1670 = _T_1669[5:0]; // @[util.scala 14:20:@231.4]
  assign _GEN_23 = _T_1670 % 6'h10; // @[util.scala 14:25:@232.4]
  assign _T_1671 = _GEN_23[4:0]; // @[util.scala 14:25:@232.4]
  assign _T_1672 = _T_1671 < _GEN_1139; // @[StoreQueue.scala 70:46:@233.4]
  assign initBits_8 = _T_1672 & io_bbStart; // @[StoreQueue.scala 70:64:@234.4]
  assign _T_1677 = 6'h19 - _GEN_1138; // @[util.scala 14:20:@236.4]
  assign _T_1678 = $unsigned(_T_1677); // @[util.scala 14:20:@237.4]
  assign _T_1679 = _T_1678[5:0]; // @[util.scala 14:20:@238.4]
  assign _GEN_24 = _T_1679 % 6'h10; // @[util.scala 14:25:@239.4]
  assign _T_1680 = _GEN_24[4:0]; // @[util.scala 14:25:@239.4]
  assign _T_1681 = _T_1680 < _GEN_1139; // @[StoreQueue.scala 70:46:@240.4]
  assign initBits_9 = _T_1681 & io_bbStart; // @[StoreQueue.scala 70:64:@241.4]
  assign _T_1686 = 6'h1a - _GEN_1138; // @[util.scala 14:20:@243.4]
  assign _T_1687 = $unsigned(_T_1686); // @[util.scala 14:20:@244.4]
  assign _T_1688 = _T_1687[5:0]; // @[util.scala 14:20:@245.4]
  assign _GEN_25 = _T_1688 % 6'h10; // @[util.scala 14:25:@246.4]
  assign _T_1689 = _GEN_25[4:0]; // @[util.scala 14:25:@246.4]
  assign _T_1690 = _T_1689 < _GEN_1139; // @[StoreQueue.scala 70:46:@247.4]
  assign initBits_10 = _T_1690 & io_bbStart; // @[StoreQueue.scala 70:64:@248.4]
  assign _T_1695 = 6'h1b - _GEN_1138; // @[util.scala 14:20:@250.4]
  assign _T_1696 = $unsigned(_T_1695); // @[util.scala 14:20:@251.4]
  assign _T_1697 = _T_1696[5:0]; // @[util.scala 14:20:@252.4]
  assign _GEN_26 = _T_1697 % 6'h10; // @[util.scala 14:25:@253.4]
  assign _T_1698 = _GEN_26[4:0]; // @[util.scala 14:25:@253.4]
  assign _T_1699 = _T_1698 < _GEN_1139; // @[StoreQueue.scala 70:46:@254.4]
  assign initBits_11 = _T_1699 & io_bbStart; // @[StoreQueue.scala 70:64:@255.4]
  assign _T_1704 = 6'h1c - _GEN_1138; // @[util.scala 14:20:@257.4]
  assign _T_1705 = $unsigned(_T_1704); // @[util.scala 14:20:@258.4]
  assign _T_1706 = _T_1705[5:0]; // @[util.scala 14:20:@259.4]
  assign _GEN_27 = _T_1706 % 6'h10; // @[util.scala 14:25:@260.4]
  assign _T_1707 = _GEN_27[4:0]; // @[util.scala 14:25:@260.4]
  assign _T_1708 = _T_1707 < _GEN_1139; // @[StoreQueue.scala 70:46:@261.4]
  assign initBits_12 = _T_1708 & io_bbStart; // @[StoreQueue.scala 70:64:@262.4]
  assign _T_1713 = 6'h1d - _GEN_1138; // @[util.scala 14:20:@264.4]
  assign _T_1714 = $unsigned(_T_1713); // @[util.scala 14:20:@265.4]
  assign _T_1715 = _T_1714[5:0]; // @[util.scala 14:20:@266.4]
  assign _GEN_28 = _T_1715 % 6'h10; // @[util.scala 14:25:@267.4]
  assign _T_1716 = _GEN_28[4:0]; // @[util.scala 14:25:@267.4]
  assign _T_1717 = _T_1716 < _GEN_1139; // @[StoreQueue.scala 70:46:@268.4]
  assign initBits_13 = _T_1717 & io_bbStart; // @[StoreQueue.scala 70:64:@269.4]
  assign _T_1722 = 6'h1e - _GEN_1138; // @[util.scala 14:20:@271.4]
  assign _T_1723 = $unsigned(_T_1722); // @[util.scala 14:20:@272.4]
  assign _T_1724 = _T_1723[5:0]; // @[util.scala 14:20:@273.4]
  assign _GEN_29 = _T_1724 % 6'h10; // @[util.scala 14:25:@274.4]
  assign _T_1725 = _GEN_29[4:0]; // @[util.scala 14:25:@274.4]
  assign _T_1726 = _T_1725 < _GEN_1139; // @[StoreQueue.scala 70:46:@275.4]
  assign initBits_14 = _T_1726 & io_bbStart; // @[StoreQueue.scala 70:64:@276.4]
  assign _T_1731 = 6'h1f - _GEN_1138; // @[util.scala 14:20:@278.4]
  assign _T_1732 = $unsigned(_T_1731); // @[util.scala 14:20:@279.4]
  assign _T_1733 = _T_1732[5:0]; // @[util.scala 14:20:@280.4]
  assign _GEN_30 = _T_1733 % 6'h10; // @[util.scala 14:25:@281.4]
  assign _T_1734 = _GEN_30[4:0]; // @[util.scala 14:25:@281.4]
  assign _T_1735 = _T_1734 < _GEN_1139; // @[StoreQueue.scala 70:46:@282.4]
  assign initBits_15 = _T_1735 & io_bbStart; // @[StoreQueue.scala 70:64:@283.4]
  assign _T_1758 = allocatedEntries_0 | initBits_0; // @[StoreQueue.scala 72:78:@301.4]
  assign _T_1759 = allocatedEntries_1 | initBits_1; // @[StoreQueue.scala 72:78:@302.4]
  assign _T_1760 = allocatedEntries_2 | initBits_2; // @[StoreQueue.scala 72:78:@303.4]
  assign _T_1761 = allocatedEntries_3 | initBits_3; // @[StoreQueue.scala 72:78:@304.4]
  assign _T_1762 = allocatedEntries_4 | initBits_4; // @[StoreQueue.scala 72:78:@305.4]
  assign _T_1763 = allocatedEntries_5 | initBits_5; // @[StoreQueue.scala 72:78:@306.4]
  assign _T_1764 = allocatedEntries_6 | initBits_6; // @[StoreQueue.scala 72:78:@307.4]
  assign _T_1765 = allocatedEntries_7 | initBits_7; // @[StoreQueue.scala 72:78:@308.4]
  assign _T_1766 = allocatedEntries_8 | initBits_8; // @[StoreQueue.scala 72:78:@309.4]
  assign _T_1767 = allocatedEntries_9 | initBits_9; // @[StoreQueue.scala 72:78:@310.4]
  assign _T_1768 = allocatedEntries_10 | initBits_10; // @[StoreQueue.scala 72:78:@311.4]
  assign _T_1769 = allocatedEntries_11 | initBits_11; // @[StoreQueue.scala 72:78:@312.4]
  assign _T_1770 = allocatedEntries_12 | initBits_12; // @[StoreQueue.scala 72:78:@313.4]
  assign _T_1771 = allocatedEntries_13 | initBits_13; // @[StoreQueue.scala 72:78:@314.4]
  assign _T_1772 = allocatedEntries_14 | initBits_14; // @[StoreQueue.scala 72:78:@315.4]
  assign _T_1773 = allocatedEntries_15 | initBits_15; // @[StoreQueue.scala 72:78:@316.4]
  assign _T_1804 = _T_1599[3:0]; // @[:@356.6]
  assign _GEN_1 = 4'h1 == _T_1804 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_2 = 4'h2 == _T_1804 ? io_bbStoreOffsets_2 : _GEN_1; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_3 = 4'h3 == _T_1804 ? io_bbStoreOffsets_3 : _GEN_2; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_4 = 4'h4 == _T_1804 ? io_bbStoreOffsets_4 : _GEN_3; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_5 = 4'h5 == _T_1804 ? io_bbStoreOffsets_5 : _GEN_4; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_6 = 4'h6 == _T_1804 ? io_bbStoreOffsets_6 : _GEN_5; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_7 = 4'h7 == _T_1804 ? io_bbStoreOffsets_7 : _GEN_6; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_8 = 4'h8 == _T_1804 ? io_bbStoreOffsets_8 : _GEN_7; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_9 = 4'h9 == _T_1804 ? io_bbStoreOffsets_9 : _GEN_8; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_10 = 4'ha == _T_1804 ? io_bbStoreOffsets_10 : _GEN_9; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_11 = 4'hb == _T_1804 ? io_bbStoreOffsets_11 : _GEN_10; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_12 = 4'hc == _T_1804 ? io_bbStoreOffsets_12 : _GEN_11; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_13 = 4'hd == _T_1804 ? io_bbStoreOffsets_13 : _GEN_12; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_14 = 4'he == _T_1804 ? io_bbStoreOffsets_14 : _GEN_13; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_15 = 4'hf == _T_1804 ? io_bbStoreOffsets_15 : _GEN_14; // @[StoreQueue.scala 76:20:@357.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[StoreQueue.scala 75:25:@350.4]
  assign _T_1822 = _T_1608[3:0]; // @[:@372.6]
  assign _GEN_35 = 4'h1 == _T_1822 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_36 = 4'h2 == _T_1822 ? io_bbStoreOffsets_2 : _GEN_35; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_37 = 4'h3 == _T_1822 ? io_bbStoreOffsets_3 : _GEN_36; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_38 = 4'h4 == _T_1822 ? io_bbStoreOffsets_4 : _GEN_37; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_39 = 4'h5 == _T_1822 ? io_bbStoreOffsets_5 : _GEN_38; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_40 = 4'h6 == _T_1822 ? io_bbStoreOffsets_6 : _GEN_39; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_41 = 4'h7 == _T_1822 ? io_bbStoreOffsets_7 : _GEN_40; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_42 = 4'h8 == _T_1822 ? io_bbStoreOffsets_8 : _GEN_41; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_43 = 4'h9 == _T_1822 ? io_bbStoreOffsets_9 : _GEN_42; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_44 = 4'ha == _T_1822 ? io_bbStoreOffsets_10 : _GEN_43; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_45 = 4'hb == _T_1822 ? io_bbStoreOffsets_11 : _GEN_44; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_46 = 4'hc == _T_1822 ? io_bbStoreOffsets_12 : _GEN_45; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_47 = 4'hd == _T_1822 ? io_bbStoreOffsets_13 : _GEN_46; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_48 = 4'he == _T_1822 ? io_bbStoreOffsets_14 : _GEN_47; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_49 = 4'hf == _T_1822 ? io_bbStoreOffsets_15 : _GEN_48; // @[StoreQueue.scala 76:20:@373.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[StoreQueue.scala 75:25:@366.4]
  assign _T_1840 = _T_1617[3:0]; // @[:@388.6]
  assign _GEN_69 = 4'h1 == _T_1840 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_70 = 4'h2 == _T_1840 ? io_bbStoreOffsets_2 : _GEN_69; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_71 = 4'h3 == _T_1840 ? io_bbStoreOffsets_3 : _GEN_70; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_72 = 4'h4 == _T_1840 ? io_bbStoreOffsets_4 : _GEN_71; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_73 = 4'h5 == _T_1840 ? io_bbStoreOffsets_5 : _GEN_72; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_74 = 4'h6 == _T_1840 ? io_bbStoreOffsets_6 : _GEN_73; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_75 = 4'h7 == _T_1840 ? io_bbStoreOffsets_7 : _GEN_74; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_76 = 4'h8 == _T_1840 ? io_bbStoreOffsets_8 : _GEN_75; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_77 = 4'h9 == _T_1840 ? io_bbStoreOffsets_9 : _GEN_76; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_78 = 4'ha == _T_1840 ? io_bbStoreOffsets_10 : _GEN_77; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_79 = 4'hb == _T_1840 ? io_bbStoreOffsets_11 : _GEN_78; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_80 = 4'hc == _T_1840 ? io_bbStoreOffsets_12 : _GEN_79; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_81 = 4'hd == _T_1840 ? io_bbStoreOffsets_13 : _GEN_80; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_82 = 4'he == _T_1840 ? io_bbStoreOffsets_14 : _GEN_81; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_83 = 4'hf == _T_1840 ? io_bbStoreOffsets_15 : _GEN_82; // @[StoreQueue.scala 76:20:@389.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[StoreQueue.scala 75:25:@382.4]
  assign _T_1858 = _T_1626[3:0]; // @[:@404.6]
  assign _GEN_103 = 4'h1 == _T_1858 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_104 = 4'h2 == _T_1858 ? io_bbStoreOffsets_2 : _GEN_103; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_105 = 4'h3 == _T_1858 ? io_bbStoreOffsets_3 : _GEN_104; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_106 = 4'h4 == _T_1858 ? io_bbStoreOffsets_4 : _GEN_105; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_107 = 4'h5 == _T_1858 ? io_bbStoreOffsets_5 : _GEN_106; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_108 = 4'h6 == _T_1858 ? io_bbStoreOffsets_6 : _GEN_107; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_109 = 4'h7 == _T_1858 ? io_bbStoreOffsets_7 : _GEN_108; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_110 = 4'h8 == _T_1858 ? io_bbStoreOffsets_8 : _GEN_109; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_111 = 4'h9 == _T_1858 ? io_bbStoreOffsets_9 : _GEN_110; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_112 = 4'ha == _T_1858 ? io_bbStoreOffsets_10 : _GEN_111; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_113 = 4'hb == _T_1858 ? io_bbStoreOffsets_11 : _GEN_112; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_114 = 4'hc == _T_1858 ? io_bbStoreOffsets_12 : _GEN_113; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_115 = 4'hd == _T_1858 ? io_bbStoreOffsets_13 : _GEN_114; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_116 = 4'he == _T_1858 ? io_bbStoreOffsets_14 : _GEN_115; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_117 = 4'hf == _T_1858 ? io_bbStoreOffsets_15 : _GEN_116; // @[StoreQueue.scala 76:20:@405.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[StoreQueue.scala 75:25:@398.4]
  assign _T_1876 = _T_1635[3:0]; // @[:@420.6]
  assign _GEN_137 = 4'h1 == _T_1876 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_138 = 4'h2 == _T_1876 ? io_bbStoreOffsets_2 : _GEN_137; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_139 = 4'h3 == _T_1876 ? io_bbStoreOffsets_3 : _GEN_138; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_140 = 4'h4 == _T_1876 ? io_bbStoreOffsets_4 : _GEN_139; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_141 = 4'h5 == _T_1876 ? io_bbStoreOffsets_5 : _GEN_140; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_142 = 4'h6 == _T_1876 ? io_bbStoreOffsets_6 : _GEN_141; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_143 = 4'h7 == _T_1876 ? io_bbStoreOffsets_7 : _GEN_142; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_144 = 4'h8 == _T_1876 ? io_bbStoreOffsets_8 : _GEN_143; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_145 = 4'h9 == _T_1876 ? io_bbStoreOffsets_9 : _GEN_144; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_146 = 4'ha == _T_1876 ? io_bbStoreOffsets_10 : _GEN_145; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_147 = 4'hb == _T_1876 ? io_bbStoreOffsets_11 : _GEN_146; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_148 = 4'hc == _T_1876 ? io_bbStoreOffsets_12 : _GEN_147; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_149 = 4'hd == _T_1876 ? io_bbStoreOffsets_13 : _GEN_148; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_150 = 4'he == _T_1876 ? io_bbStoreOffsets_14 : _GEN_149; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_151 = 4'hf == _T_1876 ? io_bbStoreOffsets_15 : _GEN_150; // @[StoreQueue.scala 76:20:@421.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[StoreQueue.scala 75:25:@414.4]
  assign _T_1894 = _T_1644[3:0]; // @[:@436.6]
  assign _GEN_171 = 4'h1 == _T_1894 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_172 = 4'h2 == _T_1894 ? io_bbStoreOffsets_2 : _GEN_171; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_173 = 4'h3 == _T_1894 ? io_bbStoreOffsets_3 : _GEN_172; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_174 = 4'h4 == _T_1894 ? io_bbStoreOffsets_4 : _GEN_173; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_175 = 4'h5 == _T_1894 ? io_bbStoreOffsets_5 : _GEN_174; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_176 = 4'h6 == _T_1894 ? io_bbStoreOffsets_6 : _GEN_175; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_177 = 4'h7 == _T_1894 ? io_bbStoreOffsets_7 : _GEN_176; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_178 = 4'h8 == _T_1894 ? io_bbStoreOffsets_8 : _GEN_177; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_179 = 4'h9 == _T_1894 ? io_bbStoreOffsets_9 : _GEN_178; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_180 = 4'ha == _T_1894 ? io_bbStoreOffsets_10 : _GEN_179; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_181 = 4'hb == _T_1894 ? io_bbStoreOffsets_11 : _GEN_180; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_182 = 4'hc == _T_1894 ? io_bbStoreOffsets_12 : _GEN_181; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_183 = 4'hd == _T_1894 ? io_bbStoreOffsets_13 : _GEN_182; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_184 = 4'he == _T_1894 ? io_bbStoreOffsets_14 : _GEN_183; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_185 = 4'hf == _T_1894 ? io_bbStoreOffsets_15 : _GEN_184; // @[StoreQueue.scala 76:20:@437.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[StoreQueue.scala 75:25:@430.4]
  assign _T_1912 = _T_1653[3:0]; // @[:@452.6]
  assign _GEN_205 = 4'h1 == _T_1912 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_206 = 4'h2 == _T_1912 ? io_bbStoreOffsets_2 : _GEN_205; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_207 = 4'h3 == _T_1912 ? io_bbStoreOffsets_3 : _GEN_206; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_208 = 4'h4 == _T_1912 ? io_bbStoreOffsets_4 : _GEN_207; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_209 = 4'h5 == _T_1912 ? io_bbStoreOffsets_5 : _GEN_208; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_210 = 4'h6 == _T_1912 ? io_bbStoreOffsets_6 : _GEN_209; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_211 = 4'h7 == _T_1912 ? io_bbStoreOffsets_7 : _GEN_210; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_212 = 4'h8 == _T_1912 ? io_bbStoreOffsets_8 : _GEN_211; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_213 = 4'h9 == _T_1912 ? io_bbStoreOffsets_9 : _GEN_212; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_214 = 4'ha == _T_1912 ? io_bbStoreOffsets_10 : _GEN_213; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_215 = 4'hb == _T_1912 ? io_bbStoreOffsets_11 : _GEN_214; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_216 = 4'hc == _T_1912 ? io_bbStoreOffsets_12 : _GEN_215; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_217 = 4'hd == _T_1912 ? io_bbStoreOffsets_13 : _GEN_216; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_218 = 4'he == _T_1912 ? io_bbStoreOffsets_14 : _GEN_217; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_219 = 4'hf == _T_1912 ? io_bbStoreOffsets_15 : _GEN_218; // @[StoreQueue.scala 76:20:@453.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[StoreQueue.scala 75:25:@446.4]
  assign _T_1930 = _T_1662[3:0]; // @[:@468.6]
  assign _GEN_239 = 4'h1 == _T_1930 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_240 = 4'h2 == _T_1930 ? io_bbStoreOffsets_2 : _GEN_239; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_241 = 4'h3 == _T_1930 ? io_bbStoreOffsets_3 : _GEN_240; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_242 = 4'h4 == _T_1930 ? io_bbStoreOffsets_4 : _GEN_241; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_243 = 4'h5 == _T_1930 ? io_bbStoreOffsets_5 : _GEN_242; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_244 = 4'h6 == _T_1930 ? io_bbStoreOffsets_6 : _GEN_243; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_245 = 4'h7 == _T_1930 ? io_bbStoreOffsets_7 : _GEN_244; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_246 = 4'h8 == _T_1930 ? io_bbStoreOffsets_8 : _GEN_245; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_247 = 4'h9 == _T_1930 ? io_bbStoreOffsets_9 : _GEN_246; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_248 = 4'ha == _T_1930 ? io_bbStoreOffsets_10 : _GEN_247; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_249 = 4'hb == _T_1930 ? io_bbStoreOffsets_11 : _GEN_248; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_250 = 4'hc == _T_1930 ? io_bbStoreOffsets_12 : _GEN_249; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_251 = 4'hd == _T_1930 ? io_bbStoreOffsets_13 : _GEN_250; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_252 = 4'he == _T_1930 ? io_bbStoreOffsets_14 : _GEN_251; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_253 = 4'hf == _T_1930 ? io_bbStoreOffsets_15 : _GEN_252; // @[StoreQueue.scala 76:20:@469.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[StoreQueue.scala 75:25:@462.4]
  assign _T_1948 = _T_1671[3:0]; // @[:@484.6]
  assign _GEN_273 = 4'h1 == _T_1948 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_274 = 4'h2 == _T_1948 ? io_bbStoreOffsets_2 : _GEN_273; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_275 = 4'h3 == _T_1948 ? io_bbStoreOffsets_3 : _GEN_274; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_276 = 4'h4 == _T_1948 ? io_bbStoreOffsets_4 : _GEN_275; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_277 = 4'h5 == _T_1948 ? io_bbStoreOffsets_5 : _GEN_276; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_278 = 4'h6 == _T_1948 ? io_bbStoreOffsets_6 : _GEN_277; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_279 = 4'h7 == _T_1948 ? io_bbStoreOffsets_7 : _GEN_278; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_280 = 4'h8 == _T_1948 ? io_bbStoreOffsets_8 : _GEN_279; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_281 = 4'h9 == _T_1948 ? io_bbStoreOffsets_9 : _GEN_280; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_282 = 4'ha == _T_1948 ? io_bbStoreOffsets_10 : _GEN_281; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_283 = 4'hb == _T_1948 ? io_bbStoreOffsets_11 : _GEN_282; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_284 = 4'hc == _T_1948 ? io_bbStoreOffsets_12 : _GEN_283; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_285 = 4'hd == _T_1948 ? io_bbStoreOffsets_13 : _GEN_284; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_286 = 4'he == _T_1948 ? io_bbStoreOffsets_14 : _GEN_285; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_287 = 4'hf == _T_1948 ? io_bbStoreOffsets_15 : _GEN_286; // @[StoreQueue.scala 76:20:@485.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[StoreQueue.scala 75:25:@478.4]
  assign _T_1966 = _T_1680[3:0]; // @[:@500.6]
  assign _GEN_307 = 4'h1 == _T_1966 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_308 = 4'h2 == _T_1966 ? io_bbStoreOffsets_2 : _GEN_307; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_309 = 4'h3 == _T_1966 ? io_bbStoreOffsets_3 : _GEN_308; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_310 = 4'h4 == _T_1966 ? io_bbStoreOffsets_4 : _GEN_309; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_311 = 4'h5 == _T_1966 ? io_bbStoreOffsets_5 : _GEN_310; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_312 = 4'h6 == _T_1966 ? io_bbStoreOffsets_6 : _GEN_311; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_313 = 4'h7 == _T_1966 ? io_bbStoreOffsets_7 : _GEN_312; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_314 = 4'h8 == _T_1966 ? io_bbStoreOffsets_8 : _GEN_313; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_315 = 4'h9 == _T_1966 ? io_bbStoreOffsets_9 : _GEN_314; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_316 = 4'ha == _T_1966 ? io_bbStoreOffsets_10 : _GEN_315; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_317 = 4'hb == _T_1966 ? io_bbStoreOffsets_11 : _GEN_316; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_318 = 4'hc == _T_1966 ? io_bbStoreOffsets_12 : _GEN_317; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_319 = 4'hd == _T_1966 ? io_bbStoreOffsets_13 : _GEN_318; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_320 = 4'he == _T_1966 ? io_bbStoreOffsets_14 : _GEN_319; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_321 = 4'hf == _T_1966 ? io_bbStoreOffsets_15 : _GEN_320; // @[StoreQueue.scala 76:20:@501.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[StoreQueue.scala 75:25:@494.4]
  assign _T_1984 = _T_1689[3:0]; // @[:@516.6]
  assign _GEN_341 = 4'h1 == _T_1984 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_342 = 4'h2 == _T_1984 ? io_bbStoreOffsets_2 : _GEN_341; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_343 = 4'h3 == _T_1984 ? io_bbStoreOffsets_3 : _GEN_342; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_344 = 4'h4 == _T_1984 ? io_bbStoreOffsets_4 : _GEN_343; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_345 = 4'h5 == _T_1984 ? io_bbStoreOffsets_5 : _GEN_344; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_346 = 4'h6 == _T_1984 ? io_bbStoreOffsets_6 : _GEN_345; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_347 = 4'h7 == _T_1984 ? io_bbStoreOffsets_7 : _GEN_346; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_348 = 4'h8 == _T_1984 ? io_bbStoreOffsets_8 : _GEN_347; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_349 = 4'h9 == _T_1984 ? io_bbStoreOffsets_9 : _GEN_348; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_350 = 4'ha == _T_1984 ? io_bbStoreOffsets_10 : _GEN_349; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_351 = 4'hb == _T_1984 ? io_bbStoreOffsets_11 : _GEN_350; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_352 = 4'hc == _T_1984 ? io_bbStoreOffsets_12 : _GEN_351; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_353 = 4'hd == _T_1984 ? io_bbStoreOffsets_13 : _GEN_352; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_354 = 4'he == _T_1984 ? io_bbStoreOffsets_14 : _GEN_353; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_355 = 4'hf == _T_1984 ? io_bbStoreOffsets_15 : _GEN_354; // @[StoreQueue.scala 76:20:@517.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[StoreQueue.scala 75:25:@510.4]
  assign _T_2002 = _T_1698[3:0]; // @[:@532.6]
  assign _GEN_375 = 4'h1 == _T_2002 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_376 = 4'h2 == _T_2002 ? io_bbStoreOffsets_2 : _GEN_375; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_377 = 4'h3 == _T_2002 ? io_bbStoreOffsets_3 : _GEN_376; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_378 = 4'h4 == _T_2002 ? io_bbStoreOffsets_4 : _GEN_377; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_379 = 4'h5 == _T_2002 ? io_bbStoreOffsets_5 : _GEN_378; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_380 = 4'h6 == _T_2002 ? io_bbStoreOffsets_6 : _GEN_379; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_381 = 4'h7 == _T_2002 ? io_bbStoreOffsets_7 : _GEN_380; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_382 = 4'h8 == _T_2002 ? io_bbStoreOffsets_8 : _GEN_381; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_383 = 4'h9 == _T_2002 ? io_bbStoreOffsets_9 : _GEN_382; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_384 = 4'ha == _T_2002 ? io_bbStoreOffsets_10 : _GEN_383; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_385 = 4'hb == _T_2002 ? io_bbStoreOffsets_11 : _GEN_384; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_386 = 4'hc == _T_2002 ? io_bbStoreOffsets_12 : _GEN_385; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_387 = 4'hd == _T_2002 ? io_bbStoreOffsets_13 : _GEN_386; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_388 = 4'he == _T_2002 ? io_bbStoreOffsets_14 : _GEN_387; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_389 = 4'hf == _T_2002 ? io_bbStoreOffsets_15 : _GEN_388; // @[StoreQueue.scala 76:20:@533.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[StoreQueue.scala 75:25:@526.4]
  assign _T_2020 = _T_1707[3:0]; // @[:@548.6]
  assign _GEN_409 = 4'h1 == _T_2020 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_410 = 4'h2 == _T_2020 ? io_bbStoreOffsets_2 : _GEN_409; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_411 = 4'h3 == _T_2020 ? io_bbStoreOffsets_3 : _GEN_410; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_412 = 4'h4 == _T_2020 ? io_bbStoreOffsets_4 : _GEN_411; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_413 = 4'h5 == _T_2020 ? io_bbStoreOffsets_5 : _GEN_412; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_414 = 4'h6 == _T_2020 ? io_bbStoreOffsets_6 : _GEN_413; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_415 = 4'h7 == _T_2020 ? io_bbStoreOffsets_7 : _GEN_414; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_416 = 4'h8 == _T_2020 ? io_bbStoreOffsets_8 : _GEN_415; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_417 = 4'h9 == _T_2020 ? io_bbStoreOffsets_9 : _GEN_416; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_418 = 4'ha == _T_2020 ? io_bbStoreOffsets_10 : _GEN_417; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_419 = 4'hb == _T_2020 ? io_bbStoreOffsets_11 : _GEN_418; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_420 = 4'hc == _T_2020 ? io_bbStoreOffsets_12 : _GEN_419; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_421 = 4'hd == _T_2020 ? io_bbStoreOffsets_13 : _GEN_420; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_422 = 4'he == _T_2020 ? io_bbStoreOffsets_14 : _GEN_421; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_423 = 4'hf == _T_2020 ? io_bbStoreOffsets_15 : _GEN_422; // @[StoreQueue.scala 76:20:@549.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[StoreQueue.scala 75:25:@542.4]
  assign _T_2038 = _T_1716[3:0]; // @[:@564.6]
  assign _GEN_443 = 4'h1 == _T_2038 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_444 = 4'h2 == _T_2038 ? io_bbStoreOffsets_2 : _GEN_443; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_445 = 4'h3 == _T_2038 ? io_bbStoreOffsets_3 : _GEN_444; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_446 = 4'h4 == _T_2038 ? io_bbStoreOffsets_4 : _GEN_445; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_447 = 4'h5 == _T_2038 ? io_bbStoreOffsets_5 : _GEN_446; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_448 = 4'h6 == _T_2038 ? io_bbStoreOffsets_6 : _GEN_447; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_449 = 4'h7 == _T_2038 ? io_bbStoreOffsets_7 : _GEN_448; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_450 = 4'h8 == _T_2038 ? io_bbStoreOffsets_8 : _GEN_449; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_451 = 4'h9 == _T_2038 ? io_bbStoreOffsets_9 : _GEN_450; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_452 = 4'ha == _T_2038 ? io_bbStoreOffsets_10 : _GEN_451; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_453 = 4'hb == _T_2038 ? io_bbStoreOffsets_11 : _GEN_452; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_454 = 4'hc == _T_2038 ? io_bbStoreOffsets_12 : _GEN_453; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_455 = 4'hd == _T_2038 ? io_bbStoreOffsets_13 : _GEN_454; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_456 = 4'he == _T_2038 ? io_bbStoreOffsets_14 : _GEN_455; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_457 = 4'hf == _T_2038 ? io_bbStoreOffsets_15 : _GEN_456; // @[StoreQueue.scala 76:20:@565.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[StoreQueue.scala 75:25:@558.4]
  assign _T_2056 = _T_1725[3:0]; // @[:@580.6]
  assign _GEN_477 = 4'h1 == _T_2056 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_478 = 4'h2 == _T_2056 ? io_bbStoreOffsets_2 : _GEN_477; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_479 = 4'h3 == _T_2056 ? io_bbStoreOffsets_3 : _GEN_478; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_480 = 4'h4 == _T_2056 ? io_bbStoreOffsets_4 : _GEN_479; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_481 = 4'h5 == _T_2056 ? io_bbStoreOffsets_5 : _GEN_480; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_482 = 4'h6 == _T_2056 ? io_bbStoreOffsets_6 : _GEN_481; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_483 = 4'h7 == _T_2056 ? io_bbStoreOffsets_7 : _GEN_482; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_484 = 4'h8 == _T_2056 ? io_bbStoreOffsets_8 : _GEN_483; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_485 = 4'h9 == _T_2056 ? io_bbStoreOffsets_9 : _GEN_484; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_486 = 4'ha == _T_2056 ? io_bbStoreOffsets_10 : _GEN_485; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_487 = 4'hb == _T_2056 ? io_bbStoreOffsets_11 : _GEN_486; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_488 = 4'hc == _T_2056 ? io_bbStoreOffsets_12 : _GEN_487; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_489 = 4'hd == _T_2056 ? io_bbStoreOffsets_13 : _GEN_488; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_490 = 4'he == _T_2056 ? io_bbStoreOffsets_14 : _GEN_489; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_491 = 4'hf == _T_2056 ? io_bbStoreOffsets_15 : _GEN_490; // @[StoreQueue.scala 76:20:@581.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[StoreQueue.scala 75:25:@574.4]
  assign _T_2074 = _T_1734[3:0]; // @[:@596.6]
  assign _GEN_511 = 4'h1 == _T_2074 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_512 = 4'h2 == _T_2074 ? io_bbStoreOffsets_2 : _GEN_511; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_513 = 4'h3 == _T_2074 ? io_bbStoreOffsets_3 : _GEN_512; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_514 = 4'h4 == _T_2074 ? io_bbStoreOffsets_4 : _GEN_513; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_515 = 4'h5 == _T_2074 ? io_bbStoreOffsets_5 : _GEN_514; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_516 = 4'h6 == _T_2074 ? io_bbStoreOffsets_6 : _GEN_515; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_517 = 4'h7 == _T_2074 ? io_bbStoreOffsets_7 : _GEN_516; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_518 = 4'h8 == _T_2074 ? io_bbStoreOffsets_8 : _GEN_517; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_519 = 4'h9 == _T_2074 ? io_bbStoreOffsets_9 : _GEN_518; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_520 = 4'ha == _T_2074 ? io_bbStoreOffsets_10 : _GEN_519; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_521 = 4'hb == _T_2074 ? io_bbStoreOffsets_11 : _GEN_520; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_522 = 4'hc == _T_2074 ? io_bbStoreOffsets_12 : _GEN_521; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_523 = 4'hd == _T_2074 ? io_bbStoreOffsets_13 : _GEN_522; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_524 = 4'he == _T_2074 ? io_bbStoreOffsets_14 : _GEN_523; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_525 = 4'hf == _T_2074 ? io_bbStoreOffsets_15 : _GEN_524; // @[StoreQueue.scala 76:20:@597.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[StoreQueue.scala 75:25:@590.4]
  assign _T_2096 = _GEN_15 + 4'h1; // @[util.scala 10:8:@615.6]
  assign _GEN_31 = _T_2096 % 5'h10; // @[util.scala 10:14:@616.6]
  assign _T_2097 = _GEN_31[4:0]; // @[util.scala 10:14:@616.6]
  assign _GEN_1203 = {{1'd0}, io_loadTail}; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2098 = _T_2097 == _GEN_1203; // @[StoreQueue.scala 96:56:@617.6]
  assign _T_2099 = io_loadEmpty & _T_2098; // @[StoreQueue.scala 95:50:@618.6]
  assign _T_2101 = _T_2099 == 1'h0; // @[StoreQueue.scala 95:35:@619.6]
  assign _T_2103 = previousLoadHead <= offsetQ_0; // @[StoreQueue.scala 100:35:@627.8]
  assign _T_2104 = offsetQ_0 < io_loadHead; // @[StoreQueue.scala 100:87:@628.8]
  assign _T_2105 = _T_2103 & _T_2104; // @[StoreQueue.scala 100:61:@629.8]
  assign _T_2107 = previousLoadHead > io_loadHead; // @[StoreQueue.scala 102:35:@634.10]
  assign _T_2108 = io_loadHead <= offsetQ_0; // @[StoreQueue.scala 103:23:@635.10]
  assign _T_2109 = offsetQ_0 < previousLoadHead; // @[StoreQueue.scala 103:75:@636.10]
  assign _T_2110 = _T_2108 & _T_2109; // @[StoreQueue.scala 103:49:@637.10]
  assign _T_2112 = _T_2110 == 1'h0; // @[StoreQueue.scala 103:9:@638.10]
  assign _T_2113 = _T_2107 & _T_2112; // @[StoreQueue.scala 102:49:@639.10]
  assign _GEN_560 = _T_2113 ? 1'h0 : checkBits_0; // @[StoreQueue.scala 103:96:@640.10]
  assign _GEN_561 = _T_2105 ? 1'h0 : _GEN_560; // @[StoreQueue.scala 100:102:@630.8]
  assign _GEN_562 = io_loadEmpty ? 1'h0 : _GEN_561; // @[StoreQueue.scala 98:26:@623.6]
  assign _GEN_563 = initBits_0 ? _T_2101 : _GEN_562; // @[StoreQueue.scala 94:35:@608.4]
  assign _T_2126 = _GEN_49 + 4'h1; // @[util.scala 10:8:@651.6]
  assign _GEN_34 = _T_2126 % 5'h10; // @[util.scala 10:14:@652.6]
  assign _T_2127 = _GEN_34[4:0]; // @[util.scala 10:14:@652.6]
  assign _T_2128 = _T_2127 == _GEN_1203; // @[StoreQueue.scala 96:56:@653.6]
  assign _T_2129 = io_loadEmpty & _T_2128; // @[StoreQueue.scala 95:50:@654.6]
  assign _T_2131 = _T_2129 == 1'h0; // @[StoreQueue.scala 95:35:@655.6]
  assign _T_2133 = previousLoadHead <= offsetQ_1; // @[StoreQueue.scala 100:35:@663.8]
  assign _T_2134 = offsetQ_1 < io_loadHead; // @[StoreQueue.scala 100:87:@664.8]
  assign _T_2135 = _T_2133 & _T_2134; // @[StoreQueue.scala 100:61:@665.8]
  assign _T_2138 = io_loadHead <= offsetQ_1; // @[StoreQueue.scala 103:23:@671.10]
  assign _T_2139 = offsetQ_1 < previousLoadHead; // @[StoreQueue.scala 103:75:@672.10]
  assign _T_2140 = _T_2138 & _T_2139; // @[StoreQueue.scala 103:49:@673.10]
  assign _T_2142 = _T_2140 == 1'h0; // @[StoreQueue.scala 103:9:@674.10]
  assign _T_2143 = _T_2107 & _T_2142; // @[StoreQueue.scala 102:49:@675.10]
  assign _GEN_580 = _T_2143 ? 1'h0 : checkBits_1; // @[StoreQueue.scala 103:96:@676.10]
  assign _GEN_581 = _T_2135 ? 1'h0 : _GEN_580; // @[StoreQueue.scala 100:102:@666.8]
  assign _GEN_582 = io_loadEmpty ? 1'h0 : _GEN_581; // @[StoreQueue.scala 98:26:@659.6]
  assign _GEN_583 = initBits_1 ? _T_2131 : _GEN_582; // @[StoreQueue.scala 94:35:@644.4]
  assign _T_2156 = _GEN_83 + 4'h1; // @[util.scala 10:8:@687.6]
  assign _GEN_50 = _T_2156 % 5'h10; // @[util.scala 10:14:@688.6]
  assign _T_2157 = _GEN_50[4:0]; // @[util.scala 10:14:@688.6]
  assign _T_2158 = _T_2157 == _GEN_1203; // @[StoreQueue.scala 96:56:@689.6]
  assign _T_2159 = io_loadEmpty & _T_2158; // @[StoreQueue.scala 95:50:@690.6]
  assign _T_2161 = _T_2159 == 1'h0; // @[StoreQueue.scala 95:35:@691.6]
  assign _T_2163 = previousLoadHead <= offsetQ_2; // @[StoreQueue.scala 100:35:@699.8]
  assign _T_2164 = offsetQ_2 < io_loadHead; // @[StoreQueue.scala 100:87:@700.8]
  assign _T_2165 = _T_2163 & _T_2164; // @[StoreQueue.scala 100:61:@701.8]
  assign _T_2168 = io_loadHead <= offsetQ_2; // @[StoreQueue.scala 103:23:@707.10]
  assign _T_2169 = offsetQ_2 < previousLoadHead; // @[StoreQueue.scala 103:75:@708.10]
  assign _T_2170 = _T_2168 & _T_2169; // @[StoreQueue.scala 103:49:@709.10]
  assign _T_2172 = _T_2170 == 1'h0; // @[StoreQueue.scala 103:9:@710.10]
  assign _T_2173 = _T_2107 & _T_2172; // @[StoreQueue.scala 102:49:@711.10]
  assign _GEN_600 = _T_2173 ? 1'h0 : checkBits_2; // @[StoreQueue.scala 103:96:@712.10]
  assign _GEN_601 = _T_2165 ? 1'h0 : _GEN_600; // @[StoreQueue.scala 100:102:@702.8]
  assign _GEN_602 = io_loadEmpty ? 1'h0 : _GEN_601; // @[StoreQueue.scala 98:26:@695.6]
  assign _GEN_603 = initBits_2 ? _T_2161 : _GEN_602; // @[StoreQueue.scala 94:35:@680.4]
  assign _T_2186 = _GEN_117 + 4'h1; // @[util.scala 10:8:@723.6]
  assign _GEN_51 = _T_2186 % 5'h10; // @[util.scala 10:14:@724.6]
  assign _T_2187 = _GEN_51[4:0]; // @[util.scala 10:14:@724.6]
  assign _T_2188 = _T_2187 == _GEN_1203; // @[StoreQueue.scala 96:56:@725.6]
  assign _T_2189 = io_loadEmpty & _T_2188; // @[StoreQueue.scala 95:50:@726.6]
  assign _T_2191 = _T_2189 == 1'h0; // @[StoreQueue.scala 95:35:@727.6]
  assign _T_2193 = previousLoadHead <= offsetQ_3; // @[StoreQueue.scala 100:35:@735.8]
  assign _T_2194 = offsetQ_3 < io_loadHead; // @[StoreQueue.scala 100:87:@736.8]
  assign _T_2195 = _T_2193 & _T_2194; // @[StoreQueue.scala 100:61:@737.8]
  assign _T_2198 = io_loadHead <= offsetQ_3; // @[StoreQueue.scala 103:23:@743.10]
  assign _T_2199 = offsetQ_3 < previousLoadHead; // @[StoreQueue.scala 103:75:@744.10]
  assign _T_2200 = _T_2198 & _T_2199; // @[StoreQueue.scala 103:49:@745.10]
  assign _T_2202 = _T_2200 == 1'h0; // @[StoreQueue.scala 103:9:@746.10]
  assign _T_2203 = _T_2107 & _T_2202; // @[StoreQueue.scala 102:49:@747.10]
  assign _GEN_620 = _T_2203 ? 1'h0 : checkBits_3; // @[StoreQueue.scala 103:96:@748.10]
  assign _GEN_621 = _T_2195 ? 1'h0 : _GEN_620; // @[StoreQueue.scala 100:102:@738.8]
  assign _GEN_622 = io_loadEmpty ? 1'h0 : _GEN_621; // @[StoreQueue.scala 98:26:@731.6]
  assign _GEN_623 = initBits_3 ? _T_2191 : _GEN_622; // @[StoreQueue.scala 94:35:@716.4]
  assign _T_2216 = _GEN_151 + 4'h1; // @[util.scala 10:8:@759.6]
  assign _GEN_52 = _T_2216 % 5'h10; // @[util.scala 10:14:@760.6]
  assign _T_2217 = _GEN_52[4:0]; // @[util.scala 10:14:@760.6]
  assign _T_2218 = _T_2217 == _GEN_1203; // @[StoreQueue.scala 96:56:@761.6]
  assign _T_2219 = io_loadEmpty & _T_2218; // @[StoreQueue.scala 95:50:@762.6]
  assign _T_2221 = _T_2219 == 1'h0; // @[StoreQueue.scala 95:35:@763.6]
  assign _T_2223 = previousLoadHead <= offsetQ_4; // @[StoreQueue.scala 100:35:@771.8]
  assign _T_2224 = offsetQ_4 < io_loadHead; // @[StoreQueue.scala 100:87:@772.8]
  assign _T_2225 = _T_2223 & _T_2224; // @[StoreQueue.scala 100:61:@773.8]
  assign _T_2228 = io_loadHead <= offsetQ_4; // @[StoreQueue.scala 103:23:@779.10]
  assign _T_2229 = offsetQ_4 < previousLoadHead; // @[StoreQueue.scala 103:75:@780.10]
  assign _T_2230 = _T_2228 & _T_2229; // @[StoreQueue.scala 103:49:@781.10]
  assign _T_2232 = _T_2230 == 1'h0; // @[StoreQueue.scala 103:9:@782.10]
  assign _T_2233 = _T_2107 & _T_2232; // @[StoreQueue.scala 102:49:@783.10]
  assign _GEN_640 = _T_2233 ? 1'h0 : checkBits_4; // @[StoreQueue.scala 103:96:@784.10]
  assign _GEN_641 = _T_2225 ? 1'h0 : _GEN_640; // @[StoreQueue.scala 100:102:@774.8]
  assign _GEN_642 = io_loadEmpty ? 1'h0 : _GEN_641; // @[StoreQueue.scala 98:26:@767.6]
  assign _GEN_643 = initBits_4 ? _T_2221 : _GEN_642; // @[StoreQueue.scala 94:35:@752.4]
  assign _T_2246 = _GEN_185 + 4'h1; // @[util.scala 10:8:@795.6]
  assign _GEN_53 = _T_2246 % 5'h10; // @[util.scala 10:14:@796.6]
  assign _T_2247 = _GEN_53[4:0]; // @[util.scala 10:14:@796.6]
  assign _T_2248 = _T_2247 == _GEN_1203; // @[StoreQueue.scala 96:56:@797.6]
  assign _T_2249 = io_loadEmpty & _T_2248; // @[StoreQueue.scala 95:50:@798.6]
  assign _T_2251 = _T_2249 == 1'h0; // @[StoreQueue.scala 95:35:@799.6]
  assign _T_2253 = previousLoadHead <= offsetQ_5; // @[StoreQueue.scala 100:35:@807.8]
  assign _T_2254 = offsetQ_5 < io_loadHead; // @[StoreQueue.scala 100:87:@808.8]
  assign _T_2255 = _T_2253 & _T_2254; // @[StoreQueue.scala 100:61:@809.8]
  assign _T_2258 = io_loadHead <= offsetQ_5; // @[StoreQueue.scala 103:23:@815.10]
  assign _T_2259 = offsetQ_5 < previousLoadHead; // @[StoreQueue.scala 103:75:@816.10]
  assign _T_2260 = _T_2258 & _T_2259; // @[StoreQueue.scala 103:49:@817.10]
  assign _T_2262 = _T_2260 == 1'h0; // @[StoreQueue.scala 103:9:@818.10]
  assign _T_2263 = _T_2107 & _T_2262; // @[StoreQueue.scala 102:49:@819.10]
  assign _GEN_660 = _T_2263 ? 1'h0 : checkBits_5; // @[StoreQueue.scala 103:96:@820.10]
  assign _GEN_661 = _T_2255 ? 1'h0 : _GEN_660; // @[StoreQueue.scala 100:102:@810.8]
  assign _GEN_662 = io_loadEmpty ? 1'h0 : _GEN_661; // @[StoreQueue.scala 98:26:@803.6]
  assign _GEN_663 = initBits_5 ? _T_2251 : _GEN_662; // @[StoreQueue.scala 94:35:@788.4]
  assign _T_2276 = _GEN_219 + 4'h1; // @[util.scala 10:8:@831.6]
  assign _GEN_54 = _T_2276 % 5'h10; // @[util.scala 10:14:@832.6]
  assign _T_2277 = _GEN_54[4:0]; // @[util.scala 10:14:@832.6]
  assign _T_2278 = _T_2277 == _GEN_1203; // @[StoreQueue.scala 96:56:@833.6]
  assign _T_2279 = io_loadEmpty & _T_2278; // @[StoreQueue.scala 95:50:@834.6]
  assign _T_2281 = _T_2279 == 1'h0; // @[StoreQueue.scala 95:35:@835.6]
  assign _T_2283 = previousLoadHead <= offsetQ_6; // @[StoreQueue.scala 100:35:@843.8]
  assign _T_2284 = offsetQ_6 < io_loadHead; // @[StoreQueue.scala 100:87:@844.8]
  assign _T_2285 = _T_2283 & _T_2284; // @[StoreQueue.scala 100:61:@845.8]
  assign _T_2288 = io_loadHead <= offsetQ_6; // @[StoreQueue.scala 103:23:@851.10]
  assign _T_2289 = offsetQ_6 < previousLoadHead; // @[StoreQueue.scala 103:75:@852.10]
  assign _T_2290 = _T_2288 & _T_2289; // @[StoreQueue.scala 103:49:@853.10]
  assign _T_2292 = _T_2290 == 1'h0; // @[StoreQueue.scala 103:9:@854.10]
  assign _T_2293 = _T_2107 & _T_2292; // @[StoreQueue.scala 102:49:@855.10]
  assign _GEN_680 = _T_2293 ? 1'h0 : checkBits_6; // @[StoreQueue.scala 103:96:@856.10]
  assign _GEN_681 = _T_2285 ? 1'h0 : _GEN_680; // @[StoreQueue.scala 100:102:@846.8]
  assign _GEN_682 = io_loadEmpty ? 1'h0 : _GEN_681; // @[StoreQueue.scala 98:26:@839.6]
  assign _GEN_683 = initBits_6 ? _T_2281 : _GEN_682; // @[StoreQueue.scala 94:35:@824.4]
  assign _T_2306 = _GEN_253 + 4'h1; // @[util.scala 10:8:@867.6]
  assign _GEN_55 = _T_2306 % 5'h10; // @[util.scala 10:14:@868.6]
  assign _T_2307 = _GEN_55[4:0]; // @[util.scala 10:14:@868.6]
  assign _T_2308 = _T_2307 == _GEN_1203; // @[StoreQueue.scala 96:56:@869.6]
  assign _T_2309 = io_loadEmpty & _T_2308; // @[StoreQueue.scala 95:50:@870.6]
  assign _T_2311 = _T_2309 == 1'h0; // @[StoreQueue.scala 95:35:@871.6]
  assign _T_2313 = previousLoadHead <= offsetQ_7; // @[StoreQueue.scala 100:35:@879.8]
  assign _T_2314 = offsetQ_7 < io_loadHead; // @[StoreQueue.scala 100:87:@880.8]
  assign _T_2315 = _T_2313 & _T_2314; // @[StoreQueue.scala 100:61:@881.8]
  assign _T_2318 = io_loadHead <= offsetQ_7; // @[StoreQueue.scala 103:23:@887.10]
  assign _T_2319 = offsetQ_7 < previousLoadHead; // @[StoreQueue.scala 103:75:@888.10]
  assign _T_2320 = _T_2318 & _T_2319; // @[StoreQueue.scala 103:49:@889.10]
  assign _T_2322 = _T_2320 == 1'h0; // @[StoreQueue.scala 103:9:@890.10]
  assign _T_2323 = _T_2107 & _T_2322; // @[StoreQueue.scala 102:49:@891.10]
  assign _GEN_700 = _T_2323 ? 1'h0 : checkBits_7; // @[StoreQueue.scala 103:96:@892.10]
  assign _GEN_701 = _T_2315 ? 1'h0 : _GEN_700; // @[StoreQueue.scala 100:102:@882.8]
  assign _GEN_702 = io_loadEmpty ? 1'h0 : _GEN_701; // @[StoreQueue.scala 98:26:@875.6]
  assign _GEN_703 = initBits_7 ? _T_2311 : _GEN_702; // @[StoreQueue.scala 94:35:@860.4]
  assign _T_2336 = _GEN_287 + 4'h1; // @[util.scala 10:8:@903.6]
  assign _GEN_56 = _T_2336 % 5'h10; // @[util.scala 10:14:@904.6]
  assign _T_2337 = _GEN_56[4:0]; // @[util.scala 10:14:@904.6]
  assign _T_2338 = _T_2337 == _GEN_1203; // @[StoreQueue.scala 96:56:@905.6]
  assign _T_2339 = io_loadEmpty & _T_2338; // @[StoreQueue.scala 95:50:@906.6]
  assign _T_2341 = _T_2339 == 1'h0; // @[StoreQueue.scala 95:35:@907.6]
  assign _T_2343 = previousLoadHead <= offsetQ_8; // @[StoreQueue.scala 100:35:@915.8]
  assign _T_2344 = offsetQ_8 < io_loadHead; // @[StoreQueue.scala 100:87:@916.8]
  assign _T_2345 = _T_2343 & _T_2344; // @[StoreQueue.scala 100:61:@917.8]
  assign _T_2348 = io_loadHead <= offsetQ_8; // @[StoreQueue.scala 103:23:@923.10]
  assign _T_2349 = offsetQ_8 < previousLoadHead; // @[StoreQueue.scala 103:75:@924.10]
  assign _T_2350 = _T_2348 & _T_2349; // @[StoreQueue.scala 103:49:@925.10]
  assign _T_2352 = _T_2350 == 1'h0; // @[StoreQueue.scala 103:9:@926.10]
  assign _T_2353 = _T_2107 & _T_2352; // @[StoreQueue.scala 102:49:@927.10]
  assign _GEN_720 = _T_2353 ? 1'h0 : checkBits_8; // @[StoreQueue.scala 103:96:@928.10]
  assign _GEN_721 = _T_2345 ? 1'h0 : _GEN_720; // @[StoreQueue.scala 100:102:@918.8]
  assign _GEN_722 = io_loadEmpty ? 1'h0 : _GEN_721; // @[StoreQueue.scala 98:26:@911.6]
  assign _GEN_723 = initBits_8 ? _T_2341 : _GEN_722; // @[StoreQueue.scala 94:35:@896.4]
  assign _T_2366 = _GEN_321 + 4'h1; // @[util.scala 10:8:@939.6]
  assign _GEN_57 = _T_2366 % 5'h10; // @[util.scala 10:14:@940.6]
  assign _T_2367 = _GEN_57[4:0]; // @[util.scala 10:14:@940.6]
  assign _T_2368 = _T_2367 == _GEN_1203; // @[StoreQueue.scala 96:56:@941.6]
  assign _T_2369 = io_loadEmpty & _T_2368; // @[StoreQueue.scala 95:50:@942.6]
  assign _T_2371 = _T_2369 == 1'h0; // @[StoreQueue.scala 95:35:@943.6]
  assign _T_2373 = previousLoadHead <= offsetQ_9; // @[StoreQueue.scala 100:35:@951.8]
  assign _T_2374 = offsetQ_9 < io_loadHead; // @[StoreQueue.scala 100:87:@952.8]
  assign _T_2375 = _T_2373 & _T_2374; // @[StoreQueue.scala 100:61:@953.8]
  assign _T_2378 = io_loadHead <= offsetQ_9; // @[StoreQueue.scala 103:23:@959.10]
  assign _T_2379 = offsetQ_9 < previousLoadHead; // @[StoreQueue.scala 103:75:@960.10]
  assign _T_2380 = _T_2378 & _T_2379; // @[StoreQueue.scala 103:49:@961.10]
  assign _T_2382 = _T_2380 == 1'h0; // @[StoreQueue.scala 103:9:@962.10]
  assign _T_2383 = _T_2107 & _T_2382; // @[StoreQueue.scala 102:49:@963.10]
  assign _GEN_740 = _T_2383 ? 1'h0 : checkBits_9; // @[StoreQueue.scala 103:96:@964.10]
  assign _GEN_741 = _T_2375 ? 1'h0 : _GEN_740; // @[StoreQueue.scala 100:102:@954.8]
  assign _GEN_742 = io_loadEmpty ? 1'h0 : _GEN_741; // @[StoreQueue.scala 98:26:@947.6]
  assign _GEN_743 = initBits_9 ? _T_2371 : _GEN_742; // @[StoreQueue.scala 94:35:@932.4]
  assign _T_2396 = _GEN_355 + 4'h1; // @[util.scala 10:8:@975.6]
  assign _GEN_58 = _T_2396 % 5'h10; // @[util.scala 10:14:@976.6]
  assign _T_2397 = _GEN_58[4:0]; // @[util.scala 10:14:@976.6]
  assign _T_2398 = _T_2397 == _GEN_1203; // @[StoreQueue.scala 96:56:@977.6]
  assign _T_2399 = io_loadEmpty & _T_2398; // @[StoreQueue.scala 95:50:@978.6]
  assign _T_2401 = _T_2399 == 1'h0; // @[StoreQueue.scala 95:35:@979.6]
  assign _T_2403 = previousLoadHead <= offsetQ_10; // @[StoreQueue.scala 100:35:@987.8]
  assign _T_2404 = offsetQ_10 < io_loadHead; // @[StoreQueue.scala 100:87:@988.8]
  assign _T_2405 = _T_2403 & _T_2404; // @[StoreQueue.scala 100:61:@989.8]
  assign _T_2408 = io_loadHead <= offsetQ_10; // @[StoreQueue.scala 103:23:@995.10]
  assign _T_2409 = offsetQ_10 < previousLoadHead; // @[StoreQueue.scala 103:75:@996.10]
  assign _T_2410 = _T_2408 & _T_2409; // @[StoreQueue.scala 103:49:@997.10]
  assign _T_2412 = _T_2410 == 1'h0; // @[StoreQueue.scala 103:9:@998.10]
  assign _T_2413 = _T_2107 & _T_2412; // @[StoreQueue.scala 102:49:@999.10]
  assign _GEN_760 = _T_2413 ? 1'h0 : checkBits_10; // @[StoreQueue.scala 103:96:@1000.10]
  assign _GEN_761 = _T_2405 ? 1'h0 : _GEN_760; // @[StoreQueue.scala 100:102:@990.8]
  assign _GEN_762 = io_loadEmpty ? 1'h0 : _GEN_761; // @[StoreQueue.scala 98:26:@983.6]
  assign _GEN_763 = initBits_10 ? _T_2401 : _GEN_762; // @[StoreQueue.scala 94:35:@968.4]
  assign _T_2426 = _GEN_389 + 4'h1; // @[util.scala 10:8:@1011.6]
  assign _GEN_59 = _T_2426 % 5'h10; // @[util.scala 10:14:@1012.6]
  assign _T_2427 = _GEN_59[4:0]; // @[util.scala 10:14:@1012.6]
  assign _T_2428 = _T_2427 == _GEN_1203; // @[StoreQueue.scala 96:56:@1013.6]
  assign _T_2429 = io_loadEmpty & _T_2428; // @[StoreQueue.scala 95:50:@1014.6]
  assign _T_2431 = _T_2429 == 1'h0; // @[StoreQueue.scala 95:35:@1015.6]
  assign _T_2433 = previousLoadHead <= offsetQ_11; // @[StoreQueue.scala 100:35:@1023.8]
  assign _T_2434 = offsetQ_11 < io_loadHead; // @[StoreQueue.scala 100:87:@1024.8]
  assign _T_2435 = _T_2433 & _T_2434; // @[StoreQueue.scala 100:61:@1025.8]
  assign _T_2438 = io_loadHead <= offsetQ_11; // @[StoreQueue.scala 103:23:@1031.10]
  assign _T_2439 = offsetQ_11 < previousLoadHead; // @[StoreQueue.scala 103:75:@1032.10]
  assign _T_2440 = _T_2438 & _T_2439; // @[StoreQueue.scala 103:49:@1033.10]
  assign _T_2442 = _T_2440 == 1'h0; // @[StoreQueue.scala 103:9:@1034.10]
  assign _T_2443 = _T_2107 & _T_2442; // @[StoreQueue.scala 102:49:@1035.10]
  assign _GEN_780 = _T_2443 ? 1'h0 : checkBits_11; // @[StoreQueue.scala 103:96:@1036.10]
  assign _GEN_781 = _T_2435 ? 1'h0 : _GEN_780; // @[StoreQueue.scala 100:102:@1026.8]
  assign _GEN_782 = io_loadEmpty ? 1'h0 : _GEN_781; // @[StoreQueue.scala 98:26:@1019.6]
  assign _GEN_783 = initBits_11 ? _T_2431 : _GEN_782; // @[StoreQueue.scala 94:35:@1004.4]
  assign _T_2456 = _GEN_423 + 4'h1; // @[util.scala 10:8:@1047.6]
  assign _GEN_60 = _T_2456 % 5'h10; // @[util.scala 10:14:@1048.6]
  assign _T_2457 = _GEN_60[4:0]; // @[util.scala 10:14:@1048.6]
  assign _T_2458 = _T_2457 == _GEN_1203; // @[StoreQueue.scala 96:56:@1049.6]
  assign _T_2459 = io_loadEmpty & _T_2458; // @[StoreQueue.scala 95:50:@1050.6]
  assign _T_2461 = _T_2459 == 1'h0; // @[StoreQueue.scala 95:35:@1051.6]
  assign _T_2463 = previousLoadHead <= offsetQ_12; // @[StoreQueue.scala 100:35:@1059.8]
  assign _T_2464 = offsetQ_12 < io_loadHead; // @[StoreQueue.scala 100:87:@1060.8]
  assign _T_2465 = _T_2463 & _T_2464; // @[StoreQueue.scala 100:61:@1061.8]
  assign _T_2468 = io_loadHead <= offsetQ_12; // @[StoreQueue.scala 103:23:@1067.10]
  assign _T_2469 = offsetQ_12 < previousLoadHead; // @[StoreQueue.scala 103:75:@1068.10]
  assign _T_2470 = _T_2468 & _T_2469; // @[StoreQueue.scala 103:49:@1069.10]
  assign _T_2472 = _T_2470 == 1'h0; // @[StoreQueue.scala 103:9:@1070.10]
  assign _T_2473 = _T_2107 & _T_2472; // @[StoreQueue.scala 102:49:@1071.10]
  assign _GEN_800 = _T_2473 ? 1'h0 : checkBits_12; // @[StoreQueue.scala 103:96:@1072.10]
  assign _GEN_801 = _T_2465 ? 1'h0 : _GEN_800; // @[StoreQueue.scala 100:102:@1062.8]
  assign _GEN_802 = io_loadEmpty ? 1'h0 : _GEN_801; // @[StoreQueue.scala 98:26:@1055.6]
  assign _GEN_803 = initBits_12 ? _T_2461 : _GEN_802; // @[StoreQueue.scala 94:35:@1040.4]
  assign _T_2486 = _GEN_457 + 4'h1; // @[util.scala 10:8:@1083.6]
  assign _GEN_61 = _T_2486 % 5'h10; // @[util.scala 10:14:@1084.6]
  assign _T_2487 = _GEN_61[4:0]; // @[util.scala 10:14:@1084.6]
  assign _T_2488 = _T_2487 == _GEN_1203; // @[StoreQueue.scala 96:56:@1085.6]
  assign _T_2489 = io_loadEmpty & _T_2488; // @[StoreQueue.scala 95:50:@1086.6]
  assign _T_2491 = _T_2489 == 1'h0; // @[StoreQueue.scala 95:35:@1087.6]
  assign _T_2493 = previousLoadHead <= offsetQ_13; // @[StoreQueue.scala 100:35:@1095.8]
  assign _T_2494 = offsetQ_13 < io_loadHead; // @[StoreQueue.scala 100:87:@1096.8]
  assign _T_2495 = _T_2493 & _T_2494; // @[StoreQueue.scala 100:61:@1097.8]
  assign _T_2498 = io_loadHead <= offsetQ_13; // @[StoreQueue.scala 103:23:@1103.10]
  assign _T_2499 = offsetQ_13 < previousLoadHead; // @[StoreQueue.scala 103:75:@1104.10]
  assign _T_2500 = _T_2498 & _T_2499; // @[StoreQueue.scala 103:49:@1105.10]
  assign _T_2502 = _T_2500 == 1'h0; // @[StoreQueue.scala 103:9:@1106.10]
  assign _T_2503 = _T_2107 & _T_2502; // @[StoreQueue.scala 102:49:@1107.10]
  assign _GEN_820 = _T_2503 ? 1'h0 : checkBits_13; // @[StoreQueue.scala 103:96:@1108.10]
  assign _GEN_821 = _T_2495 ? 1'h0 : _GEN_820; // @[StoreQueue.scala 100:102:@1098.8]
  assign _GEN_822 = io_loadEmpty ? 1'h0 : _GEN_821; // @[StoreQueue.scala 98:26:@1091.6]
  assign _GEN_823 = initBits_13 ? _T_2491 : _GEN_822; // @[StoreQueue.scala 94:35:@1076.4]
  assign _T_2516 = _GEN_491 + 4'h1; // @[util.scala 10:8:@1119.6]
  assign _GEN_62 = _T_2516 % 5'h10; // @[util.scala 10:14:@1120.6]
  assign _T_2517 = _GEN_62[4:0]; // @[util.scala 10:14:@1120.6]
  assign _T_2518 = _T_2517 == _GEN_1203; // @[StoreQueue.scala 96:56:@1121.6]
  assign _T_2519 = io_loadEmpty & _T_2518; // @[StoreQueue.scala 95:50:@1122.6]
  assign _T_2521 = _T_2519 == 1'h0; // @[StoreQueue.scala 95:35:@1123.6]
  assign _T_2523 = previousLoadHead <= offsetQ_14; // @[StoreQueue.scala 100:35:@1131.8]
  assign _T_2524 = offsetQ_14 < io_loadHead; // @[StoreQueue.scala 100:87:@1132.8]
  assign _T_2525 = _T_2523 & _T_2524; // @[StoreQueue.scala 100:61:@1133.8]
  assign _T_2528 = io_loadHead <= offsetQ_14; // @[StoreQueue.scala 103:23:@1139.10]
  assign _T_2529 = offsetQ_14 < previousLoadHead; // @[StoreQueue.scala 103:75:@1140.10]
  assign _T_2530 = _T_2528 & _T_2529; // @[StoreQueue.scala 103:49:@1141.10]
  assign _T_2532 = _T_2530 == 1'h0; // @[StoreQueue.scala 103:9:@1142.10]
  assign _T_2533 = _T_2107 & _T_2532; // @[StoreQueue.scala 102:49:@1143.10]
  assign _GEN_840 = _T_2533 ? 1'h0 : checkBits_14; // @[StoreQueue.scala 103:96:@1144.10]
  assign _GEN_841 = _T_2525 ? 1'h0 : _GEN_840; // @[StoreQueue.scala 100:102:@1134.8]
  assign _GEN_842 = io_loadEmpty ? 1'h0 : _GEN_841; // @[StoreQueue.scala 98:26:@1127.6]
  assign _GEN_843 = initBits_14 ? _T_2521 : _GEN_842; // @[StoreQueue.scala 94:35:@1112.4]
  assign _T_2546 = _GEN_525 + 4'h1; // @[util.scala 10:8:@1155.6]
  assign _GEN_63 = _T_2546 % 5'h10; // @[util.scala 10:14:@1156.6]
  assign _T_2547 = _GEN_63[4:0]; // @[util.scala 10:14:@1156.6]
  assign _T_2548 = _T_2547 == _GEN_1203; // @[StoreQueue.scala 96:56:@1157.6]
  assign _T_2549 = io_loadEmpty & _T_2548; // @[StoreQueue.scala 95:50:@1158.6]
  assign _T_2551 = _T_2549 == 1'h0; // @[StoreQueue.scala 95:35:@1159.6]
  assign _T_2553 = previousLoadHead <= offsetQ_15; // @[StoreQueue.scala 100:35:@1167.8]
  assign _T_2554 = offsetQ_15 < io_loadHead; // @[StoreQueue.scala 100:87:@1168.8]
  assign _T_2555 = _T_2553 & _T_2554; // @[StoreQueue.scala 100:61:@1169.8]
  assign _T_2558 = io_loadHead <= offsetQ_15; // @[StoreQueue.scala 103:23:@1175.10]
  assign _T_2559 = offsetQ_15 < previousLoadHead; // @[StoreQueue.scala 103:75:@1176.10]
  assign _T_2560 = _T_2558 & _T_2559; // @[StoreQueue.scala 103:49:@1177.10]
  assign _T_2562 = _T_2560 == 1'h0; // @[StoreQueue.scala 103:9:@1178.10]
  assign _T_2563 = _T_2107 & _T_2562; // @[StoreQueue.scala 102:49:@1179.10]
  assign _GEN_860 = _T_2563 ? 1'h0 : checkBits_15; // @[StoreQueue.scala 103:96:@1180.10]
  assign _GEN_861 = _T_2555 ? 1'h0 : _GEN_860; // @[StoreQueue.scala 100:102:@1170.8]
  assign _GEN_862 = io_loadEmpty ? 1'h0 : _GEN_861; // @[StoreQueue.scala 98:26:@1163.6]
  assign _GEN_863 = initBits_15 ? _T_2551 : _GEN_862; // @[StoreQueue.scala 94:35:@1148.4]
  assign _T_2565 = io_loadHead < io_loadTail; // @[StoreQueue.scala 119:103:@1184.4]
  assign _T_2567 = io_loadHead <= 4'h0; // @[StoreQueue.scala 120:17:@1185.4]
  assign _T_2569 = 4'h0 < io_loadTail; // @[StoreQueue.scala 120:35:@1186.4]
  assign _T_2570 = _T_2567 & _T_2569; // @[StoreQueue.scala 120:26:@1187.4]
  assign _T_2572 = io_loadEmpty == 1'h0; // @[StoreQueue.scala 120:50:@1188.4]
  assign _T_2574 = io_loadTail <= 4'h0; // @[StoreQueue.scala 120:81:@1189.4]
  assign _T_2576 = 4'h0 < io_loadHead; // @[StoreQueue.scala 120:99:@1190.4]
  assign _T_2577 = _T_2574 & _T_2576; // @[StoreQueue.scala 120:90:@1191.4]
  assign _T_2579 = _T_2577 == 1'h0; // @[StoreQueue.scala 120:67:@1192.4]
  assign _T_2580 = _T_2572 & _T_2579; // @[StoreQueue.scala 120:64:@1193.4]
  assign validEntriesInLoadQ_0 = _T_2565 ? _T_2570 : _T_2580; // @[StoreQueue.scala 119:90:@1194.4]
  assign _T_2584 = io_loadHead <= 4'h1; // @[StoreQueue.scala 120:17:@1196.4]
  assign _T_2586 = 4'h1 < io_loadTail; // @[StoreQueue.scala 120:35:@1197.4]
  assign _T_2587 = _T_2584 & _T_2586; // @[StoreQueue.scala 120:26:@1198.4]
  assign _T_2591 = io_loadTail <= 4'h1; // @[StoreQueue.scala 120:81:@1200.4]
  assign _T_2593 = 4'h1 < io_loadHead; // @[StoreQueue.scala 120:99:@1201.4]
  assign _T_2594 = _T_2591 & _T_2593; // @[StoreQueue.scala 120:90:@1202.4]
  assign _T_2596 = _T_2594 == 1'h0; // @[StoreQueue.scala 120:67:@1203.4]
  assign _T_2597 = _T_2572 & _T_2596; // @[StoreQueue.scala 120:64:@1204.4]
  assign validEntriesInLoadQ_1 = _T_2565 ? _T_2587 : _T_2597; // @[StoreQueue.scala 119:90:@1205.4]
  assign _T_2601 = io_loadHead <= 4'h2; // @[StoreQueue.scala 120:17:@1207.4]
  assign _T_2603 = 4'h2 < io_loadTail; // @[StoreQueue.scala 120:35:@1208.4]
  assign _T_2604 = _T_2601 & _T_2603; // @[StoreQueue.scala 120:26:@1209.4]
  assign _T_2608 = io_loadTail <= 4'h2; // @[StoreQueue.scala 120:81:@1211.4]
  assign _T_2610 = 4'h2 < io_loadHead; // @[StoreQueue.scala 120:99:@1212.4]
  assign _T_2611 = _T_2608 & _T_2610; // @[StoreQueue.scala 120:90:@1213.4]
  assign _T_2613 = _T_2611 == 1'h0; // @[StoreQueue.scala 120:67:@1214.4]
  assign _T_2614 = _T_2572 & _T_2613; // @[StoreQueue.scala 120:64:@1215.4]
  assign validEntriesInLoadQ_2 = _T_2565 ? _T_2604 : _T_2614; // @[StoreQueue.scala 119:90:@1216.4]
  assign _T_2618 = io_loadHead <= 4'h3; // @[StoreQueue.scala 120:17:@1218.4]
  assign _T_2620 = 4'h3 < io_loadTail; // @[StoreQueue.scala 120:35:@1219.4]
  assign _T_2621 = _T_2618 & _T_2620; // @[StoreQueue.scala 120:26:@1220.4]
  assign _T_2625 = io_loadTail <= 4'h3; // @[StoreQueue.scala 120:81:@1222.4]
  assign _T_2627 = 4'h3 < io_loadHead; // @[StoreQueue.scala 120:99:@1223.4]
  assign _T_2628 = _T_2625 & _T_2627; // @[StoreQueue.scala 120:90:@1224.4]
  assign _T_2630 = _T_2628 == 1'h0; // @[StoreQueue.scala 120:67:@1225.4]
  assign _T_2631 = _T_2572 & _T_2630; // @[StoreQueue.scala 120:64:@1226.4]
  assign validEntriesInLoadQ_3 = _T_2565 ? _T_2621 : _T_2631; // @[StoreQueue.scala 119:90:@1227.4]
  assign _T_2635 = io_loadHead <= 4'h4; // @[StoreQueue.scala 120:17:@1229.4]
  assign _T_2637 = 4'h4 < io_loadTail; // @[StoreQueue.scala 120:35:@1230.4]
  assign _T_2638 = _T_2635 & _T_2637; // @[StoreQueue.scala 120:26:@1231.4]
  assign _T_2642 = io_loadTail <= 4'h4; // @[StoreQueue.scala 120:81:@1233.4]
  assign _T_2644 = 4'h4 < io_loadHead; // @[StoreQueue.scala 120:99:@1234.4]
  assign _T_2645 = _T_2642 & _T_2644; // @[StoreQueue.scala 120:90:@1235.4]
  assign _T_2647 = _T_2645 == 1'h0; // @[StoreQueue.scala 120:67:@1236.4]
  assign _T_2648 = _T_2572 & _T_2647; // @[StoreQueue.scala 120:64:@1237.4]
  assign validEntriesInLoadQ_4 = _T_2565 ? _T_2638 : _T_2648; // @[StoreQueue.scala 119:90:@1238.4]
  assign _T_2652 = io_loadHead <= 4'h5; // @[StoreQueue.scala 120:17:@1240.4]
  assign _T_2654 = 4'h5 < io_loadTail; // @[StoreQueue.scala 120:35:@1241.4]
  assign _T_2655 = _T_2652 & _T_2654; // @[StoreQueue.scala 120:26:@1242.4]
  assign _T_2659 = io_loadTail <= 4'h5; // @[StoreQueue.scala 120:81:@1244.4]
  assign _T_2661 = 4'h5 < io_loadHead; // @[StoreQueue.scala 120:99:@1245.4]
  assign _T_2662 = _T_2659 & _T_2661; // @[StoreQueue.scala 120:90:@1246.4]
  assign _T_2664 = _T_2662 == 1'h0; // @[StoreQueue.scala 120:67:@1247.4]
  assign _T_2665 = _T_2572 & _T_2664; // @[StoreQueue.scala 120:64:@1248.4]
  assign validEntriesInLoadQ_5 = _T_2565 ? _T_2655 : _T_2665; // @[StoreQueue.scala 119:90:@1249.4]
  assign _T_2669 = io_loadHead <= 4'h6; // @[StoreQueue.scala 120:17:@1251.4]
  assign _T_2671 = 4'h6 < io_loadTail; // @[StoreQueue.scala 120:35:@1252.4]
  assign _T_2672 = _T_2669 & _T_2671; // @[StoreQueue.scala 120:26:@1253.4]
  assign _T_2676 = io_loadTail <= 4'h6; // @[StoreQueue.scala 120:81:@1255.4]
  assign _T_2678 = 4'h6 < io_loadHead; // @[StoreQueue.scala 120:99:@1256.4]
  assign _T_2679 = _T_2676 & _T_2678; // @[StoreQueue.scala 120:90:@1257.4]
  assign _T_2681 = _T_2679 == 1'h0; // @[StoreQueue.scala 120:67:@1258.4]
  assign _T_2682 = _T_2572 & _T_2681; // @[StoreQueue.scala 120:64:@1259.4]
  assign validEntriesInLoadQ_6 = _T_2565 ? _T_2672 : _T_2682; // @[StoreQueue.scala 119:90:@1260.4]
  assign _T_2686 = io_loadHead <= 4'h7; // @[StoreQueue.scala 120:17:@1262.4]
  assign _T_2688 = 4'h7 < io_loadTail; // @[StoreQueue.scala 120:35:@1263.4]
  assign _T_2689 = _T_2686 & _T_2688; // @[StoreQueue.scala 120:26:@1264.4]
  assign _T_2693 = io_loadTail <= 4'h7; // @[StoreQueue.scala 120:81:@1266.4]
  assign _T_2695 = 4'h7 < io_loadHead; // @[StoreQueue.scala 120:99:@1267.4]
  assign _T_2696 = _T_2693 & _T_2695; // @[StoreQueue.scala 120:90:@1268.4]
  assign _T_2698 = _T_2696 == 1'h0; // @[StoreQueue.scala 120:67:@1269.4]
  assign _T_2699 = _T_2572 & _T_2698; // @[StoreQueue.scala 120:64:@1270.4]
  assign validEntriesInLoadQ_7 = _T_2565 ? _T_2689 : _T_2699; // @[StoreQueue.scala 119:90:@1271.4]
  assign _T_2703 = io_loadHead <= 4'h8; // @[StoreQueue.scala 120:17:@1273.4]
  assign _T_2705 = 4'h8 < io_loadTail; // @[StoreQueue.scala 120:35:@1274.4]
  assign _T_2706 = _T_2703 & _T_2705; // @[StoreQueue.scala 120:26:@1275.4]
  assign _T_2710 = io_loadTail <= 4'h8; // @[StoreQueue.scala 120:81:@1277.4]
  assign _T_2712 = 4'h8 < io_loadHead; // @[StoreQueue.scala 120:99:@1278.4]
  assign _T_2713 = _T_2710 & _T_2712; // @[StoreQueue.scala 120:90:@1279.4]
  assign _T_2715 = _T_2713 == 1'h0; // @[StoreQueue.scala 120:67:@1280.4]
  assign _T_2716 = _T_2572 & _T_2715; // @[StoreQueue.scala 120:64:@1281.4]
  assign validEntriesInLoadQ_8 = _T_2565 ? _T_2706 : _T_2716; // @[StoreQueue.scala 119:90:@1282.4]
  assign _T_2720 = io_loadHead <= 4'h9; // @[StoreQueue.scala 120:17:@1284.4]
  assign _T_2722 = 4'h9 < io_loadTail; // @[StoreQueue.scala 120:35:@1285.4]
  assign _T_2723 = _T_2720 & _T_2722; // @[StoreQueue.scala 120:26:@1286.4]
  assign _T_2727 = io_loadTail <= 4'h9; // @[StoreQueue.scala 120:81:@1288.4]
  assign _T_2729 = 4'h9 < io_loadHead; // @[StoreQueue.scala 120:99:@1289.4]
  assign _T_2730 = _T_2727 & _T_2729; // @[StoreQueue.scala 120:90:@1290.4]
  assign _T_2732 = _T_2730 == 1'h0; // @[StoreQueue.scala 120:67:@1291.4]
  assign _T_2733 = _T_2572 & _T_2732; // @[StoreQueue.scala 120:64:@1292.4]
  assign validEntriesInLoadQ_9 = _T_2565 ? _T_2723 : _T_2733; // @[StoreQueue.scala 119:90:@1293.4]
  assign _T_2737 = io_loadHead <= 4'ha; // @[StoreQueue.scala 120:17:@1295.4]
  assign _T_2739 = 4'ha < io_loadTail; // @[StoreQueue.scala 120:35:@1296.4]
  assign _T_2740 = _T_2737 & _T_2739; // @[StoreQueue.scala 120:26:@1297.4]
  assign _T_2744 = io_loadTail <= 4'ha; // @[StoreQueue.scala 120:81:@1299.4]
  assign _T_2746 = 4'ha < io_loadHead; // @[StoreQueue.scala 120:99:@1300.4]
  assign _T_2747 = _T_2744 & _T_2746; // @[StoreQueue.scala 120:90:@1301.4]
  assign _T_2749 = _T_2747 == 1'h0; // @[StoreQueue.scala 120:67:@1302.4]
  assign _T_2750 = _T_2572 & _T_2749; // @[StoreQueue.scala 120:64:@1303.4]
  assign validEntriesInLoadQ_10 = _T_2565 ? _T_2740 : _T_2750; // @[StoreQueue.scala 119:90:@1304.4]
  assign _T_2754 = io_loadHead <= 4'hb; // @[StoreQueue.scala 120:17:@1306.4]
  assign _T_2756 = 4'hb < io_loadTail; // @[StoreQueue.scala 120:35:@1307.4]
  assign _T_2757 = _T_2754 & _T_2756; // @[StoreQueue.scala 120:26:@1308.4]
  assign _T_2761 = io_loadTail <= 4'hb; // @[StoreQueue.scala 120:81:@1310.4]
  assign _T_2763 = 4'hb < io_loadHead; // @[StoreQueue.scala 120:99:@1311.4]
  assign _T_2764 = _T_2761 & _T_2763; // @[StoreQueue.scala 120:90:@1312.4]
  assign _T_2766 = _T_2764 == 1'h0; // @[StoreQueue.scala 120:67:@1313.4]
  assign _T_2767 = _T_2572 & _T_2766; // @[StoreQueue.scala 120:64:@1314.4]
  assign validEntriesInLoadQ_11 = _T_2565 ? _T_2757 : _T_2767; // @[StoreQueue.scala 119:90:@1315.4]
  assign _T_2771 = io_loadHead <= 4'hc; // @[StoreQueue.scala 120:17:@1317.4]
  assign _T_2773 = 4'hc < io_loadTail; // @[StoreQueue.scala 120:35:@1318.4]
  assign _T_2774 = _T_2771 & _T_2773; // @[StoreQueue.scala 120:26:@1319.4]
  assign _T_2778 = io_loadTail <= 4'hc; // @[StoreQueue.scala 120:81:@1321.4]
  assign _T_2780 = 4'hc < io_loadHead; // @[StoreQueue.scala 120:99:@1322.4]
  assign _T_2781 = _T_2778 & _T_2780; // @[StoreQueue.scala 120:90:@1323.4]
  assign _T_2783 = _T_2781 == 1'h0; // @[StoreQueue.scala 120:67:@1324.4]
  assign _T_2784 = _T_2572 & _T_2783; // @[StoreQueue.scala 120:64:@1325.4]
  assign validEntriesInLoadQ_12 = _T_2565 ? _T_2774 : _T_2784; // @[StoreQueue.scala 119:90:@1326.4]
  assign _T_2788 = io_loadHead <= 4'hd; // @[StoreQueue.scala 120:17:@1328.4]
  assign _T_2790 = 4'hd < io_loadTail; // @[StoreQueue.scala 120:35:@1329.4]
  assign _T_2791 = _T_2788 & _T_2790; // @[StoreQueue.scala 120:26:@1330.4]
  assign _T_2795 = io_loadTail <= 4'hd; // @[StoreQueue.scala 120:81:@1332.4]
  assign _T_2797 = 4'hd < io_loadHead; // @[StoreQueue.scala 120:99:@1333.4]
  assign _T_2798 = _T_2795 & _T_2797; // @[StoreQueue.scala 120:90:@1334.4]
  assign _T_2800 = _T_2798 == 1'h0; // @[StoreQueue.scala 120:67:@1335.4]
  assign _T_2801 = _T_2572 & _T_2800; // @[StoreQueue.scala 120:64:@1336.4]
  assign validEntriesInLoadQ_13 = _T_2565 ? _T_2791 : _T_2801; // @[StoreQueue.scala 119:90:@1337.4]
  assign _T_2805 = io_loadHead <= 4'he; // @[StoreQueue.scala 120:17:@1339.4]
  assign _T_2807 = 4'he < io_loadTail; // @[StoreQueue.scala 120:35:@1340.4]
  assign _T_2808 = _T_2805 & _T_2807; // @[StoreQueue.scala 120:26:@1341.4]
  assign _T_2812 = io_loadTail <= 4'he; // @[StoreQueue.scala 120:81:@1343.4]
  assign _T_2814 = 4'he < io_loadHead; // @[StoreQueue.scala 120:99:@1344.4]
  assign _T_2815 = _T_2812 & _T_2814; // @[StoreQueue.scala 120:90:@1345.4]
  assign _T_2817 = _T_2815 == 1'h0; // @[StoreQueue.scala 120:67:@1346.4]
  assign _T_2818 = _T_2572 & _T_2817; // @[StoreQueue.scala 120:64:@1347.4]
  assign validEntriesInLoadQ_14 = _T_2565 ? _T_2808 : _T_2818; // @[StoreQueue.scala 119:90:@1348.4]
  assign validEntriesInLoadQ_15 = _T_2565 ? 1'h0 : _T_2572; // @[StoreQueue.scala 119:90:@1359.4]
  assign _GEN_865 = 4'h1 == head ? offsetQ_1 : offsetQ_0; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_866 = 4'h2 == head ? offsetQ_2 : _GEN_865; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_867 = 4'h3 == head ? offsetQ_3 : _GEN_866; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_868 = 4'h4 == head ? offsetQ_4 : _GEN_867; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_869 = 4'h5 == head ? offsetQ_5 : _GEN_868; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_870 = 4'h6 == head ? offsetQ_6 : _GEN_869; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_871 = 4'h7 == head ? offsetQ_7 : _GEN_870; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_872 = 4'h8 == head ? offsetQ_8 : _GEN_871; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_873 = 4'h9 == head ? offsetQ_9 : _GEN_872; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_874 = 4'ha == head ? offsetQ_10 : _GEN_873; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_875 = 4'hb == head ? offsetQ_11 : _GEN_874; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_876 = 4'hc == head ? offsetQ_12 : _GEN_875; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_877 = 4'hd == head ? offsetQ_13 : _GEN_876; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_878 = 4'he == head ? offsetQ_14 : _GEN_877; // @[StoreQueue.scala 126:96:@1377.4]
  assign _GEN_879 = 4'hf == head ? offsetQ_15 : _GEN_878; // @[StoreQueue.scala 126:96:@1377.4]
  assign _T_2861 = io_loadHead <= _GEN_879; // @[StoreQueue.scala 126:96:@1377.4]
  assign loadsToCheck_0 = _T_2861 ? _T_2567 : 1'h1; // @[StoreQueue.scala 126:83:@1385.4]
  assign _T_2891 = 4'h1 <= _GEN_879; // @[StoreQueue.scala 127:37:@1388.4]
  assign _T_2892 = _T_2584 & _T_2891; // @[StoreQueue.scala 127:28:@1389.4]
  assign _T_2897 = _GEN_879 < 4'h1; // @[StoreQueue.scala 127:71:@1390.4]
  assign _T_2900 = _T_2897 & _T_2593; // @[StoreQueue.scala 127:79:@1392.4]
  assign _T_2902 = _T_2900 == 1'h0; // @[StoreQueue.scala 127:55:@1393.4]
  assign loadsToCheck_1 = _T_2861 ? _T_2892 : _T_2902; // @[StoreQueue.scala 126:83:@1394.4]
  assign _T_2914 = 4'h2 <= _GEN_879; // @[StoreQueue.scala 127:37:@1397.4]
  assign _T_2915 = _T_2601 & _T_2914; // @[StoreQueue.scala 127:28:@1398.4]
  assign _T_2920 = _GEN_879 < 4'h2; // @[StoreQueue.scala 127:71:@1399.4]
  assign _T_2923 = _T_2920 & _T_2610; // @[StoreQueue.scala 127:79:@1401.4]
  assign _T_2925 = _T_2923 == 1'h0; // @[StoreQueue.scala 127:55:@1402.4]
  assign loadsToCheck_2 = _T_2861 ? _T_2915 : _T_2925; // @[StoreQueue.scala 126:83:@1403.4]
  assign _T_2937 = 4'h3 <= _GEN_879; // @[StoreQueue.scala 127:37:@1406.4]
  assign _T_2938 = _T_2618 & _T_2937; // @[StoreQueue.scala 127:28:@1407.4]
  assign _T_2943 = _GEN_879 < 4'h3; // @[StoreQueue.scala 127:71:@1408.4]
  assign _T_2946 = _T_2943 & _T_2627; // @[StoreQueue.scala 127:79:@1410.4]
  assign _T_2948 = _T_2946 == 1'h0; // @[StoreQueue.scala 127:55:@1411.4]
  assign loadsToCheck_3 = _T_2861 ? _T_2938 : _T_2948; // @[StoreQueue.scala 126:83:@1412.4]
  assign _T_2960 = 4'h4 <= _GEN_879; // @[StoreQueue.scala 127:37:@1415.4]
  assign _T_2961 = _T_2635 & _T_2960; // @[StoreQueue.scala 127:28:@1416.4]
  assign _T_2966 = _GEN_879 < 4'h4; // @[StoreQueue.scala 127:71:@1417.4]
  assign _T_2969 = _T_2966 & _T_2644; // @[StoreQueue.scala 127:79:@1419.4]
  assign _T_2971 = _T_2969 == 1'h0; // @[StoreQueue.scala 127:55:@1420.4]
  assign loadsToCheck_4 = _T_2861 ? _T_2961 : _T_2971; // @[StoreQueue.scala 126:83:@1421.4]
  assign _T_2983 = 4'h5 <= _GEN_879; // @[StoreQueue.scala 127:37:@1424.4]
  assign _T_2984 = _T_2652 & _T_2983; // @[StoreQueue.scala 127:28:@1425.4]
  assign _T_2989 = _GEN_879 < 4'h5; // @[StoreQueue.scala 127:71:@1426.4]
  assign _T_2992 = _T_2989 & _T_2661; // @[StoreQueue.scala 127:79:@1428.4]
  assign _T_2994 = _T_2992 == 1'h0; // @[StoreQueue.scala 127:55:@1429.4]
  assign loadsToCheck_5 = _T_2861 ? _T_2984 : _T_2994; // @[StoreQueue.scala 126:83:@1430.4]
  assign _T_3006 = 4'h6 <= _GEN_879; // @[StoreQueue.scala 127:37:@1433.4]
  assign _T_3007 = _T_2669 & _T_3006; // @[StoreQueue.scala 127:28:@1434.4]
  assign _T_3012 = _GEN_879 < 4'h6; // @[StoreQueue.scala 127:71:@1435.4]
  assign _T_3015 = _T_3012 & _T_2678; // @[StoreQueue.scala 127:79:@1437.4]
  assign _T_3017 = _T_3015 == 1'h0; // @[StoreQueue.scala 127:55:@1438.4]
  assign loadsToCheck_6 = _T_2861 ? _T_3007 : _T_3017; // @[StoreQueue.scala 126:83:@1439.4]
  assign _T_3029 = 4'h7 <= _GEN_879; // @[StoreQueue.scala 127:37:@1442.4]
  assign _T_3030 = _T_2686 & _T_3029; // @[StoreQueue.scala 127:28:@1443.4]
  assign _T_3035 = _GEN_879 < 4'h7; // @[StoreQueue.scala 127:71:@1444.4]
  assign _T_3038 = _T_3035 & _T_2695; // @[StoreQueue.scala 127:79:@1446.4]
  assign _T_3040 = _T_3038 == 1'h0; // @[StoreQueue.scala 127:55:@1447.4]
  assign loadsToCheck_7 = _T_2861 ? _T_3030 : _T_3040; // @[StoreQueue.scala 126:83:@1448.4]
  assign _T_3052 = 4'h8 <= _GEN_879; // @[StoreQueue.scala 127:37:@1451.4]
  assign _T_3053 = _T_2703 & _T_3052; // @[StoreQueue.scala 127:28:@1452.4]
  assign _T_3058 = _GEN_879 < 4'h8; // @[StoreQueue.scala 127:71:@1453.4]
  assign _T_3061 = _T_3058 & _T_2712; // @[StoreQueue.scala 127:79:@1455.4]
  assign _T_3063 = _T_3061 == 1'h0; // @[StoreQueue.scala 127:55:@1456.4]
  assign loadsToCheck_8 = _T_2861 ? _T_3053 : _T_3063; // @[StoreQueue.scala 126:83:@1457.4]
  assign _T_3075 = 4'h9 <= _GEN_879; // @[StoreQueue.scala 127:37:@1460.4]
  assign _T_3076 = _T_2720 & _T_3075; // @[StoreQueue.scala 127:28:@1461.4]
  assign _T_3081 = _GEN_879 < 4'h9; // @[StoreQueue.scala 127:71:@1462.4]
  assign _T_3084 = _T_3081 & _T_2729; // @[StoreQueue.scala 127:79:@1464.4]
  assign _T_3086 = _T_3084 == 1'h0; // @[StoreQueue.scala 127:55:@1465.4]
  assign loadsToCheck_9 = _T_2861 ? _T_3076 : _T_3086; // @[StoreQueue.scala 126:83:@1466.4]
  assign _T_3098 = 4'ha <= _GEN_879; // @[StoreQueue.scala 127:37:@1469.4]
  assign _T_3099 = _T_2737 & _T_3098; // @[StoreQueue.scala 127:28:@1470.4]
  assign _T_3104 = _GEN_879 < 4'ha; // @[StoreQueue.scala 127:71:@1471.4]
  assign _T_3107 = _T_3104 & _T_2746; // @[StoreQueue.scala 127:79:@1473.4]
  assign _T_3109 = _T_3107 == 1'h0; // @[StoreQueue.scala 127:55:@1474.4]
  assign loadsToCheck_10 = _T_2861 ? _T_3099 : _T_3109; // @[StoreQueue.scala 126:83:@1475.4]
  assign _T_3121 = 4'hb <= _GEN_879; // @[StoreQueue.scala 127:37:@1478.4]
  assign _T_3122 = _T_2754 & _T_3121; // @[StoreQueue.scala 127:28:@1479.4]
  assign _T_3127 = _GEN_879 < 4'hb; // @[StoreQueue.scala 127:71:@1480.4]
  assign _T_3130 = _T_3127 & _T_2763; // @[StoreQueue.scala 127:79:@1482.4]
  assign _T_3132 = _T_3130 == 1'h0; // @[StoreQueue.scala 127:55:@1483.4]
  assign loadsToCheck_11 = _T_2861 ? _T_3122 : _T_3132; // @[StoreQueue.scala 126:83:@1484.4]
  assign _T_3144 = 4'hc <= _GEN_879; // @[StoreQueue.scala 127:37:@1487.4]
  assign _T_3145 = _T_2771 & _T_3144; // @[StoreQueue.scala 127:28:@1488.4]
  assign _T_3150 = _GEN_879 < 4'hc; // @[StoreQueue.scala 127:71:@1489.4]
  assign _T_3153 = _T_3150 & _T_2780; // @[StoreQueue.scala 127:79:@1491.4]
  assign _T_3155 = _T_3153 == 1'h0; // @[StoreQueue.scala 127:55:@1492.4]
  assign loadsToCheck_12 = _T_2861 ? _T_3145 : _T_3155; // @[StoreQueue.scala 126:83:@1493.4]
  assign _T_3167 = 4'hd <= _GEN_879; // @[StoreQueue.scala 127:37:@1496.4]
  assign _T_3168 = _T_2788 & _T_3167; // @[StoreQueue.scala 127:28:@1497.4]
  assign _T_3173 = _GEN_879 < 4'hd; // @[StoreQueue.scala 127:71:@1498.4]
  assign _T_3176 = _T_3173 & _T_2797; // @[StoreQueue.scala 127:79:@1500.4]
  assign _T_3178 = _T_3176 == 1'h0; // @[StoreQueue.scala 127:55:@1501.4]
  assign loadsToCheck_13 = _T_2861 ? _T_3168 : _T_3178; // @[StoreQueue.scala 126:83:@1502.4]
  assign _T_3190 = 4'he <= _GEN_879; // @[StoreQueue.scala 127:37:@1505.4]
  assign _T_3191 = _T_2805 & _T_3190; // @[StoreQueue.scala 127:28:@1506.4]
  assign _T_3196 = _GEN_879 < 4'he; // @[StoreQueue.scala 127:71:@1507.4]
  assign _T_3199 = _T_3196 & _T_2814; // @[StoreQueue.scala 127:79:@1509.4]
  assign _T_3201 = _T_3199 == 1'h0; // @[StoreQueue.scala 127:55:@1510.4]
  assign loadsToCheck_14 = _T_2861 ? _T_3191 : _T_3201; // @[StoreQueue.scala 126:83:@1511.4]
  assign _T_3213 = 4'hf <= _GEN_879; // @[StoreQueue.scala 127:37:@1514.4]
  assign loadsToCheck_15 = _T_2861 ? _T_3213 : 1'h1; // @[StoreQueue.scala 126:83:@1520.4]
  assign _T_3247 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[StoreQueue.scala 133:16:@1538.4]
  assign _GEN_881 = 4'h1 == head ? checkBits_1 : checkBits_0; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_882 = 4'h2 == head ? checkBits_2 : _GEN_881; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_883 = 4'h3 == head ? checkBits_3 : _GEN_882; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_884 = 4'h4 == head ? checkBits_4 : _GEN_883; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_885 = 4'h5 == head ? checkBits_5 : _GEN_884; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_886 = 4'h6 == head ? checkBits_6 : _GEN_885; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_887 = 4'h7 == head ? checkBits_7 : _GEN_886; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_888 = 4'h8 == head ? checkBits_8 : _GEN_887; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_889 = 4'h9 == head ? checkBits_9 : _GEN_888; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_890 = 4'ha == head ? checkBits_10 : _GEN_889; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_891 = 4'hb == head ? checkBits_11 : _GEN_890; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_892 = 4'hc == head ? checkBits_12 : _GEN_891; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_893 = 4'hd == head ? checkBits_13 : _GEN_892; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_894 = 4'he == head ? checkBits_14 : _GEN_893; // @[StoreQueue.scala 133:24:@1539.4]
  assign _GEN_895 = 4'hf == head ? checkBits_15 : _GEN_894; // @[StoreQueue.scala 133:24:@1539.4]
  assign entriesToCheck_0 = _T_3247 & _GEN_895; // @[StoreQueue.scala 133:24:@1539.4]
  assign _T_3252 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[StoreQueue.scala 133:16:@1540.4]
  assign entriesToCheck_1 = _T_3252 & _GEN_895; // @[StoreQueue.scala 133:24:@1541.4]
  assign _T_3257 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[StoreQueue.scala 133:16:@1542.4]
  assign entriesToCheck_2 = _T_3257 & _GEN_895; // @[StoreQueue.scala 133:24:@1543.4]
  assign _T_3262 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[StoreQueue.scala 133:16:@1544.4]
  assign entriesToCheck_3 = _T_3262 & _GEN_895; // @[StoreQueue.scala 133:24:@1545.4]
  assign _T_3267 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[StoreQueue.scala 133:16:@1546.4]
  assign entriesToCheck_4 = _T_3267 & _GEN_895; // @[StoreQueue.scala 133:24:@1547.4]
  assign _T_3272 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[StoreQueue.scala 133:16:@1548.4]
  assign entriesToCheck_5 = _T_3272 & _GEN_895; // @[StoreQueue.scala 133:24:@1549.4]
  assign _T_3277 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[StoreQueue.scala 133:16:@1550.4]
  assign entriesToCheck_6 = _T_3277 & _GEN_895; // @[StoreQueue.scala 133:24:@1551.4]
  assign _T_3282 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[StoreQueue.scala 133:16:@1552.4]
  assign entriesToCheck_7 = _T_3282 & _GEN_895; // @[StoreQueue.scala 133:24:@1553.4]
  assign _T_3287 = loadsToCheck_8 & validEntriesInLoadQ_8; // @[StoreQueue.scala 133:16:@1554.4]
  assign entriesToCheck_8 = _T_3287 & _GEN_895; // @[StoreQueue.scala 133:24:@1555.4]
  assign _T_3292 = loadsToCheck_9 & validEntriesInLoadQ_9; // @[StoreQueue.scala 133:16:@1556.4]
  assign entriesToCheck_9 = _T_3292 & _GEN_895; // @[StoreQueue.scala 133:24:@1557.4]
  assign _T_3297 = loadsToCheck_10 & validEntriesInLoadQ_10; // @[StoreQueue.scala 133:16:@1558.4]
  assign entriesToCheck_10 = _T_3297 & _GEN_895; // @[StoreQueue.scala 133:24:@1559.4]
  assign _T_3302 = loadsToCheck_11 & validEntriesInLoadQ_11; // @[StoreQueue.scala 133:16:@1560.4]
  assign entriesToCheck_11 = _T_3302 & _GEN_895; // @[StoreQueue.scala 133:24:@1561.4]
  assign _T_3307 = loadsToCheck_12 & validEntriesInLoadQ_12; // @[StoreQueue.scala 133:16:@1562.4]
  assign entriesToCheck_12 = _T_3307 & _GEN_895; // @[StoreQueue.scala 133:24:@1563.4]
  assign _T_3312 = loadsToCheck_13 & validEntriesInLoadQ_13; // @[StoreQueue.scala 133:16:@1564.4]
  assign entriesToCheck_13 = _T_3312 & _GEN_895; // @[StoreQueue.scala 133:24:@1565.4]
  assign _T_3317 = loadsToCheck_14 & validEntriesInLoadQ_14; // @[StoreQueue.scala 133:16:@1566.4]
  assign entriesToCheck_14 = _T_3317 & _GEN_895; // @[StoreQueue.scala 133:24:@1567.4]
  assign _T_3322 = loadsToCheck_15 & validEntriesInLoadQ_15; // @[StoreQueue.scala 133:16:@1568.4]
  assign entriesToCheck_15 = _T_3322 & _GEN_895; // @[StoreQueue.scala 133:24:@1569.4]
  assign _T_3370 = entriesToCheck_0 == 1'h0; // @[StoreQueue.scala 140:34:@1588.4]
  assign _T_3371 = _T_3370 | io_loadDataDone_0; // @[StoreQueue.scala 140:64:@1589.4]
  assign _GEN_897 = 4'h1 == head ? addrQ_1 : addrQ_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_898 = 4'h2 == head ? addrQ_2 : _GEN_897; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_899 = 4'h3 == head ? addrQ_3 : _GEN_898; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_900 = 4'h4 == head ? addrQ_4 : _GEN_899; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_901 = 4'h5 == head ? addrQ_5 : _GEN_900; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_902 = 4'h6 == head ? addrQ_6 : _GEN_901; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_903 = 4'h7 == head ? addrQ_7 : _GEN_902; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_904 = 4'h8 == head ? addrQ_8 : _GEN_903; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_905 = 4'h9 == head ? addrQ_9 : _GEN_904; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_906 = 4'ha == head ? addrQ_10 : _GEN_905; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_907 = 4'hb == head ? addrQ_11 : _GEN_906; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_908 = 4'hc == head ? addrQ_12 : _GEN_907; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_909 = 4'hd == head ? addrQ_13 : _GEN_908; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_910 = 4'he == head ? addrQ_14 : _GEN_909; // @[StoreQueue.scala 141:51:@1590.4]
  assign _GEN_911 = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3375 = _GEN_911 != io_loadAddressQueue_0; // @[StoreQueue.scala 141:51:@1590.4]
  assign _T_3376 = io_loadAddressDone_0 & _T_3375; // @[StoreQueue.scala 141:36:@1591.4]
  assign noConflicts_0 = _T_3371 | _T_3376; // @[StoreQueue.scala 140:95:@1592.4]
  assign _T_3379 = entriesToCheck_1 == 1'h0; // @[StoreQueue.scala 140:34:@1594.4]
  assign _T_3380 = _T_3379 | io_loadDataDone_1; // @[StoreQueue.scala 140:64:@1595.4]
  assign _T_3384 = _GEN_911 != io_loadAddressQueue_1; // @[StoreQueue.scala 141:51:@1596.4]
  assign _T_3385 = io_loadAddressDone_1 & _T_3384; // @[StoreQueue.scala 141:36:@1597.4]
  assign noConflicts_1 = _T_3380 | _T_3385; // @[StoreQueue.scala 140:95:@1598.4]
  assign _T_3388 = entriesToCheck_2 == 1'h0; // @[StoreQueue.scala 140:34:@1600.4]
  assign _T_3389 = _T_3388 | io_loadDataDone_2; // @[StoreQueue.scala 140:64:@1601.4]
  assign _T_3393 = _GEN_911 != io_loadAddressQueue_2; // @[StoreQueue.scala 141:51:@1602.4]
  assign _T_3394 = io_loadAddressDone_2 & _T_3393; // @[StoreQueue.scala 141:36:@1603.4]
  assign noConflicts_2 = _T_3389 | _T_3394; // @[StoreQueue.scala 140:95:@1604.4]
  assign _T_3397 = entriesToCheck_3 == 1'h0; // @[StoreQueue.scala 140:34:@1606.4]
  assign _T_3398 = _T_3397 | io_loadDataDone_3; // @[StoreQueue.scala 140:64:@1607.4]
  assign _T_3402 = _GEN_911 != io_loadAddressQueue_3; // @[StoreQueue.scala 141:51:@1608.4]
  assign _T_3403 = io_loadAddressDone_3 & _T_3402; // @[StoreQueue.scala 141:36:@1609.4]
  assign noConflicts_3 = _T_3398 | _T_3403; // @[StoreQueue.scala 140:95:@1610.4]
  assign _T_3406 = entriesToCheck_4 == 1'h0; // @[StoreQueue.scala 140:34:@1612.4]
  assign _T_3407 = _T_3406 | io_loadDataDone_4; // @[StoreQueue.scala 140:64:@1613.4]
  assign _T_3411 = _GEN_911 != io_loadAddressQueue_4; // @[StoreQueue.scala 141:51:@1614.4]
  assign _T_3412 = io_loadAddressDone_4 & _T_3411; // @[StoreQueue.scala 141:36:@1615.4]
  assign noConflicts_4 = _T_3407 | _T_3412; // @[StoreQueue.scala 140:95:@1616.4]
  assign _T_3415 = entriesToCheck_5 == 1'h0; // @[StoreQueue.scala 140:34:@1618.4]
  assign _T_3416 = _T_3415 | io_loadDataDone_5; // @[StoreQueue.scala 140:64:@1619.4]
  assign _T_3420 = _GEN_911 != io_loadAddressQueue_5; // @[StoreQueue.scala 141:51:@1620.4]
  assign _T_3421 = io_loadAddressDone_5 & _T_3420; // @[StoreQueue.scala 141:36:@1621.4]
  assign noConflicts_5 = _T_3416 | _T_3421; // @[StoreQueue.scala 140:95:@1622.4]
  assign _T_3424 = entriesToCheck_6 == 1'h0; // @[StoreQueue.scala 140:34:@1624.4]
  assign _T_3425 = _T_3424 | io_loadDataDone_6; // @[StoreQueue.scala 140:64:@1625.4]
  assign _T_3429 = _GEN_911 != io_loadAddressQueue_6; // @[StoreQueue.scala 141:51:@1626.4]
  assign _T_3430 = io_loadAddressDone_6 & _T_3429; // @[StoreQueue.scala 141:36:@1627.4]
  assign noConflicts_6 = _T_3425 | _T_3430; // @[StoreQueue.scala 140:95:@1628.4]
  assign _T_3433 = entriesToCheck_7 == 1'h0; // @[StoreQueue.scala 140:34:@1630.4]
  assign _T_3434 = _T_3433 | io_loadDataDone_7; // @[StoreQueue.scala 140:64:@1631.4]
  assign _T_3438 = _GEN_911 != io_loadAddressQueue_7; // @[StoreQueue.scala 141:51:@1632.4]
  assign _T_3439 = io_loadAddressDone_7 & _T_3438; // @[StoreQueue.scala 141:36:@1633.4]
  assign noConflicts_7 = _T_3434 | _T_3439; // @[StoreQueue.scala 140:95:@1634.4]
  assign _T_3442 = entriesToCheck_8 == 1'h0; // @[StoreQueue.scala 140:34:@1636.4]
  assign _T_3443 = _T_3442 | io_loadDataDone_8; // @[StoreQueue.scala 140:64:@1637.4]
  assign _T_3447 = _GEN_911 != io_loadAddressQueue_8; // @[StoreQueue.scala 141:51:@1638.4]
  assign _T_3448 = io_loadAddressDone_8 & _T_3447; // @[StoreQueue.scala 141:36:@1639.4]
  assign noConflicts_8 = _T_3443 | _T_3448; // @[StoreQueue.scala 140:95:@1640.4]
  assign _T_3451 = entriesToCheck_9 == 1'h0; // @[StoreQueue.scala 140:34:@1642.4]
  assign _T_3452 = _T_3451 | io_loadDataDone_9; // @[StoreQueue.scala 140:64:@1643.4]
  assign _T_3456 = _GEN_911 != io_loadAddressQueue_9; // @[StoreQueue.scala 141:51:@1644.4]
  assign _T_3457 = io_loadAddressDone_9 & _T_3456; // @[StoreQueue.scala 141:36:@1645.4]
  assign noConflicts_9 = _T_3452 | _T_3457; // @[StoreQueue.scala 140:95:@1646.4]
  assign _T_3460 = entriesToCheck_10 == 1'h0; // @[StoreQueue.scala 140:34:@1648.4]
  assign _T_3461 = _T_3460 | io_loadDataDone_10; // @[StoreQueue.scala 140:64:@1649.4]
  assign _T_3465 = _GEN_911 != io_loadAddressQueue_10; // @[StoreQueue.scala 141:51:@1650.4]
  assign _T_3466 = io_loadAddressDone_10 & _T_3465; // @[StoreQueue.scala 141:36:@1651.4]
  assign noConflicts_10 = _T_3461 | _T_3466; // @[StoreQueue.scala 140:95:@1652.4]
  assign _T_3469 = entriesToCheck_11 == 1'h0; // @[StoreQueue.scala 140:34:@1654.4]
  assign _T_3470 = _T_3469 | io_loadDataDone_11; // @[StoreQueue.scala 140:64:@1655.4]
  assign _T_3474 = _GEN_911 != io_loadAddressQueue_11; // @[StoreQueue.scala 141:51:@1656.4]
  assign _T_3475 = io_loadAddressDone_11 & _T_3474; // @[StoreQueue.scala 141:36:@1657.4]
  assign noConflicts_11 = _T_3470 | _T_3475; // @[StoreQueue.scala 140:95:@1658.4]
  assign _T_3478 = entriesToCheck_12 == 1'h0; // @[StoreQueue.scala 140:34:@1660.4]
  assign _T_3479 = _T_3478 | io_loadDataDone_12; // @[StoreQueue.scala 140:64:@1661.4]
  assign _T_3483 = _GEN_911 != io_loadAddressQueue_12; // @[StoreQueue.scala 141:51:@1662.4]
  assign _T_3484 = io_loadAddressDone_12 & _T_3483; // @[StoreQueue.scala 141:36:@1663.4]
  assign noConflicts_12 = _T_3479 | _T_3484; // @[StoreQueue.scala 140:95:@1664.4]
  assign _T_3487 = entriesToCheck_13 == 1'h0; // @[StoreQueue.scala 140:34:@1666.4]
  assign _T_3488 = _T_3487 | io_loadDataDone_13; // @[StoreQueue.scala 140:64:@1667.4]
  assign _T_3492 = _GEN_911 != io_loadAddressQueue_13; // @[StoreQueue.scala 141:51:@1668.4]
  assign _T_3493 = io_loadAddressDone_13 & _T_3492; // @[StoreQueue.scala 141:36:@1669.4]
  assign noConflicts_13 = _T_3488 | _T_3493; // @[StoreQueue.scala 140:95:@1670.4]
  assign _T_3496 = entriesToCheck_14 == 1'h0; // @[StoreQueue.scala 140:34:@1672.4]
  assign _T_3497 = _T_3496 | io_loadDataDone_14; // @[StoreQueue.scala 140:64:@1673.4]
  assign _T_3501 = _GEN_911 != io_loadAddressQueue_14; // @[StoreQueue.scala 141:51:@1674.4]
  assign _T_3502 = io_loadAddressDone_14 & _T_3501; // @[StoreQueue.scala 141:36:@1675.4]
  assign noConflicts_14 = _T_3497 | _T_3502; // @[StoreQueue.scala 140:95:@1676.4]
  assign _T_3505 = entriesToCheck_15 == 1'h0; // @[StoreQueue.scala 140:34:@1678.4]
  assign _T_3506 = _T_3505 | io_loadDataDone_15; // @[StoreQueue.scala 140:64:@1679.4]
  assign _T_3510 = _GEN_911 != io_loadAddressQueue_15; // @[StoreQueue.scala 141:51:@1680.4]
  assign _T_3511 = io_loadAddressDone_15 & _T_3510; // @[StoreQueue.scala 141:36:@1681.4]
  assign noConflicts_15 = _T_3506 | _T_3511; // @[StoreQueue.scala 140:95:@1682.4]
  assign _GEN_913 = 4'h1 == head ? addrKnown_1 : addrKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_914 = 4'h2 == head ? addrKnown_2 : _GEN_913; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_915 = 4'h3 == head ? addrKnown_3 : _GEN_914; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_916 = 4'h4 == head ? addrKnown_4 : _GEN_915; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_917 = 4'h5 == head ? addrKnown_5 : _GEN_916; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_918 = 4'h6 == head ? addrKnown_6 : _GEN_917; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_919 = 4'h7 == head ? addrKnown_7 : _GEN_918; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_920 = 4'h8 == head ? addrKnown_8 : _GEN_919; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_921 = 4'h9 == head ? addrKnown_9 : _GEN_920; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_922 = 4'ha == head ? addrKnown_10 : _GEN_921; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_923 = 4'hb == head ? addrKnown_11 : _GEN_922; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_924 = 4'hc == head ? addrKnown_12 : _GEN_923; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_925 = 4'hd == head ? addrKnown_13 : _GEN_924; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_926 = 4'he == head ? addrKnown_14 : _GEN_925; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_927 = 4'hf == head ? addrKnown_15 : _GEN_926; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_929 = 4'h1 == head ? dataKnown_1 : dataKnown_0; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_930 = 4'h2 == head ? dataKnown_2 : _GEN_929; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_931 = 4'h3 == head ? dataKnown_3 : _GEN_930; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_932 = 4'h4 == head ? dataKnown_4 : _GEN_931; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_933 = 4'h5 == head ? dataKnown_5 : _GEN_932; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_934 = 4'h6 == head ? dataKnown_6 : _GEN_933; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_935 = 4'h7 == head ? dataKnown_7 : _GEN_934; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_936 = 4'h8 == head ? dataKnown_8 : _GEN_935; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_937 = 4'h9 == head ? dataKnown_9 : _GEN_936; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_938 = 4'ha == head ? dataKnown_10 : _GEN_937; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_939 = 4'hb == head ? dataKnown_11 : _GEN_938; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_940 = 4'hc == head ? dataKnown_12 : _GEN_939; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_941 = 4'hd == head ? dataKnown_13 : _GEN_940; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_942 = 4'he == head ? dataKnown_14 : _GEN_941; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_943 = 4'hf == head ? dataKnown_15 : _GEN_942; // @[StoreQueue.scala 154:44:@1684.4]
  assign _T_3519 = _GEN_927 & _GEN_943; // @[StoreQueue.scala 154:44:@1684.4]
  assign _GEN_945 = 4'h1 == head ? storeCompleted_1 : storeCompleted_0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_946 = 4'h2 == head ? storeCompleted_2 : _GEN_945; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_947 = 4'h3 == head ? storeCompleted_3 : _GEN_946; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_948 = 4'h4 == head ? storeCompleted_4 : _GEN_947; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_949 = 4'h5 == head ? storeCompleted_5 : _GEN_948; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_950 = 4'h6 == head ? storeCompleted_6 : _GEN_949; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_951 = 4'h7 == head ? storeCompleted_7 : _GEN_950; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_952 = 4'h8 == head ? storeCompleted_8 : _GEN_951; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_953 = 4'h9 == head ? storeCompleted_9 : _GEN_952; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_954 = 4'ha == head ? storeCompleted_10 : _GEN_953; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_955 = 4'hb == head ? storeCompleted_11 : _GEN_954; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_956 = 4'hc == head ? storeCompleted_12 : _GEN_955; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_957 = 4'hd == head ? storeCompleted_13 : _GEN_956; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_958 = 4'he == head ? storeCompleted_14 : _GEN_957; // @[StoreQueue.scala 154:66:@1685.4]
  assign _GEN_959 = 4'hf == head ? storeCompleted_15 : _GEN_958; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3524 = _GEN_959 == 1'h0; // @[StoreQueue.scala 154:66:@1685.4]
  assign _T_3525 = _T_3519 & _T_3524; // @[StoreQueue.scala 154:63:@1686.4]
  assign _T_3528 = noConflicts_0 & noConflicts_1; // @[StoreQueue.scala 154:109:@1688.4]
  assign _T_3529 = _T_3528 & noConflicts_2; // @[StoreQueue.scala 154:109:@1689.4]
  assign _T_3530 = _T_3529 & noConflicts_3; // @[StoreQueue.scala 154:109:@1690.4]
  assign _T_3531 = _T_3530 & noConflicts_4; // @[StoreQueue.scala 154:109:@1691.4]
  assign _T_3532 = _T_3531 & noConflicts_5; // @[StoreQueue.scala 154:109:@1692.4]
  assign _T_3533 = _T_3532 & noConflicts_6; // @[StoreQueue.scala 154:109:@1693.4]
  assign _T_3534 = _T_3533 & noConflicts_7; // @[StoreQueue.scala 154:109:@1694.4]
  assign _T_3535 = _T_3534 & noConflicts_8; // @[StoreQueue.scala 154:109:@1695.4]
  assign _T_3536 = _T_3535 & noConflicts_9; // @[StoreQueue.scala 154:109:@1696.4]
  assign _T_3537 = _T_3536 & noConflicts_10; // @[StoreQueue.scala 154:109:@1697.4]
  assign _T_3538 = _T_3537 & noConflicts_11; // @[StoreQueue.scala 154:109:@1698.4]
  assign _T_3539 = _T_3538 & noConflicts_12; // @[StoreQueue.scala 154:109:@1699.4]
  assign _T_3540 = _T_3539 & noConflicts_13; // @[StoreQueue.scala 154:109:@1700.4]
  assign _T_3541 = _T_3540 & noConflicts_14; // @[StoreQueue.scala 154:109:@1701.4]
  assign _T_3542 = _T_3541 & noConflicts_15; // @[StoreQueue.scala 154:109:@1702.4]
  assign storeRequest = _T_3525 & _T_3542; // @[StoreQueue.scala 154:88:@1703.4]
  assign _T_3545 = head == 4'h0; // @[StoreQueue.scala 164:23:@1708.6]
  assign _T_3546 = _T_3545 & storeRequest; // @[StoreQueue.scala 164:43:@1709.6]
  assign _T_3547 = _T_3546 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1710.6]
  assign _GEN_960 = _T_3547 ? 1'h1 : storeCompleted_0; // @[StoreQueue.scala 164:86:@1711.6]
  assign _GEN_961 = initBits_0 ? 1'h0 : _GEN_960; // @[StoreQueue.scala 162:37:@1704.4]
  assign _T_3551 = head == 4'h1; // @[StoreQueue.scala 164:23:@1718.6]
  assign _T_3552 = _T_3551 & storeRequest; // @[StoreQueue.scala 164:43:@1719.6]
  assign _T_3553 = _T_3552 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1720.6]
  assign _GEN_962 = _T_3553 ? 1'h1 : storeCompleted_1; // @[StoreQueue.scala 164:86:@1721.6]
  assign _GEN_963 = initBits_1 ? 1'h0 : _GEN_962; // @[StoreQueue.scala 162:37:@1714.4]
  assign _T_3557 = head == 4'h2; // @[StoreQueue.scala 164:23:@1728.6]
  assign _T_3558 = _T_3557 & storeRequest; // @[StoreQueue.scala 164:43:@1729.6]
  assign _T_3559 = _T_3558 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1730.6]
  assign _GEN_964 = _T_3559 ? 1'h1 : storeCompleted_2; // @[StoreQueue.scala 164:86:@1731.6]
  assign _GEN_965 = initBits_2 ? 1'h0 : _GEN_964; // @[StoreQueue.scala 162:37:@1724.4]
  assign _T_3563 = head == 4'h3; // @[StoreQueue.scala 164:23:@1738.6]
  assign _T_3564 = _T_3563 & storeRequest; // @[StoreQueue.scala 164:43:@1739.6]
  assign _T_3565 = _T_3564 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1740.6]
  assign _GEN_966 = _T_3565 ? 1'h1 : storeCompleted_3; // @[StoreQueue.scala 164:86:@1741.6]
  assign _GEN_967 = initBits_3 ? 1'h0 : _GEN_966; // @[StoreQueue.scala 162:37:@1734.4]
  assign _T_3569 = head == 4'h4; // @[StoreQueue.scala 164:23:@1748.6]
  assign _T_3570 = _T_3569 & storeRequest; // @[StoreQueue.scala 164:43:@1749.6]
  assign _T_3571 = _T_3570 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1750.6]
  assign _GEN_968 = _T_3571 ? 1'h1 : storeCompleted_4; // @[StoreQueue.scala 164:86:@1751.6]
  assign _GEN_969 = initBits_4 ? 1'h0 : _GEN_968; // @[StoreQueue.scala 162:37:@1744.4]
  assign _T_3575 = head == 4'h5; // @[StoreQueue.scala 164:23:@1758.6]
  assign _T_3576 = _T_3575 & storeRequest; // @[StoreQueue.scala 164:43:@1759.6]
  assign _T_3577 = _T_3576 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1760.6]
  assign _GEN_970 = _T_3577 ? 1'h1 : storeCompleted_5; // @[StoreQueue.scala 164:86:@1761.6]
  assign _GEN_971 = initBits_5 ? 1'h0 : _GEN_970; // @[StoreQueue.scala 162:37:@1754.4]
  assign _T_3581 = head == 4'h6; // @[StoreQueue.scala 164:23:@1768.6]
  assign _T_3582 = _T_3581 & storeRequest; // @[StoreQueue.scala 164:43:@1769.6]
  assign _T_3583 = _T_3582 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1770.6]
  assign _GEN_972 = _T_3583 ? 1'h1 : storeCompleted_6; // @[StoreQueue.scala 164:86:@1771.6]
  assign _GEN_973 = initBits_6 ? 1'h0 : _GEN_972; // @[StoreQueue.scala 162:37:@1764.4]
  assign _T_3587 = head == 4'h7; // @[StoreQueue.scala 164:23:@1778.6]
  assign _T_3588 = _T_3587 & storeRequest; // @[StoreQueue.scala 164:43:@1779.6]
  assign _T_3589 = _T_3588 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1780.6]
  assign _GEN_974 = _T_3589 ? 1'h1 : storeCompleted_7; // @[StoreQueue.scala 164:86:@1781.6]
  assign _GEN_975 = initBits_7 ? 1'h0 : _GEN_974; // @[StoreQueue.scala 162:37:@1774.4]
  assign _T_3593 = head == 4'h8; // @[StoreQueue.scala 164:23:@1788.6]
  assign _T_3594 = _T_3593 & storeRequest; // @[StoreQueue.scala 164:43:@1789.6]
  assign _T_3595 = _T_3594 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1790.6]
  assign _GEN_976 = _T_3595 ? 1'h1 : storeCompleted_8; // @[StoreQueue.scala 164:86:@1791.6]
  assign _GEN_977 = initBits_8 ? 1'h0 : _GEN_976; // @[StoreQueue.scala 162:37:@1784.4]
  assign _T_3599 = head == 4'h9; // @[StoreQueue.scala 164:23:@1798.6]
  assign _T_3600 = _T_3599 & storeRequest; // @[StoreQueue.scala 164:43:@1799.6]
  assign _T_3601 = _T_3600 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1800.6]
  assign _GEN_978 = _T_3601 ? 1'h1 : storeCompleted_9; // @[StoreQueue.scala 164:86:@1801.6]
  assign _GEN_979 = initBits_9 ? 1'h0 : _GEN_978; // @[StoreQueue.scala 162:37:@1794.4]
  assign _T_3605 = head == 4'ha; // @[StoreQueue.scala 164:23:@1808.6]
  assign _T_3606 = _T_3605 & storeRequest; // @[StoreQueue.scala 164:43:@1809.6]
  assign _T_3607 = _T_3606 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1810.6]
  assign _GEN_980 = _T_3607 ? 1'h1 : storeCompleted_10; // @[StoreQueue.scala 164:86:@1811.6]
  assign _GEN_981 = initBits_10 ? 1'h0 : _GEN_980; // @[StoreQueue.scala 162:37:@1804.4]
  assign _T_3611 = head == 4'hb; // @[StoreQueue.scala 164:23:@1818.6]
  assign _T_3612 = _T_3611 & storeRequest; // @[StoreQueue.scala 164:43:@1819.6]
  assign _T_3613 = _T_3612 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1820.6]
  assign _GEN_982 = _T_3613 ? 1'h1 : storeCompleted_11; // @[StoreQueue.scala 164:86:@1821.6]
  assign _GEN_983 = initBits_11 ? 1'h0 : _GEN_982; // @[StoreQueue.scala 162:37:@1814.4]
  assign _T_3617 = head == 4'hc; // @[StoreQueue.scala 164:23:@1828.6]
  assign _T_3618 = _T_3617 & storeRequest; // @[StoreQueue.scala 164:43:@1829.6]
  assign _T_3619 = _T_3618 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1830.6]
  assign _GEN_984 = _T_3619 ? 1'h1 : storeCompleted_12; // @[StoreQueue.scala 164:86:@1831.6]
  assign _GEN_985 = initBits_12 ? 1'h0 : _GEN_984; // @[StoreQueue.scala 162:37:@1824.4]
  assign _T_3623 = head == 4'hd; // @[StoreQueue.scala 164:23:@1838.6]
  assign _T_3624 = _T_3623 & storeRequest; // @[StoreQueue.scala 164:43:@1839.6]
  assign _T_3625 = _T_3624 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1840.6]
  assign _GEN_986 = _T_3625 ? 1'h1 : storeCompleted_13; // @[StoreQueue.scala 164:86:@1841.6]
  assign _GEN_987 = initBits_13 ? 1'h0 : _GEN_986; // @[StoreQueue.scala 162:37:@1834.4]
  assign _T_3629 = head == 4'he; // @[StoreQueue.scala 164:23:@1848.6]
  assign _T_3630 = _T_3629 & storeRequest; // @[StoreQueue.scala 164:43:@1849.6]
  assign _T_3631 = _T_3630 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1850.6]
  assign _GEN_988 = _T_3631 ? 1'h1 : storeCompleted_14; // @[StoreQueue.scala 164:86:@1851.6]
  assign _GEN_989 = initBits_14 ? 1'h0 : _GEN_988; // @[StoreQueue.scala 162:37:@1844.4]
  assign _T_3635 = head == 4'hf; // @[StoreQueue.scala 164:23:@1858.6]
  assign _T_3636 = _T_3635 & storeRequest; // @[StoreQueue.scala 164:43:@1859.6]
  assign _T_3637 = _T_3636 & io_memIsReadyForStores; // @[StoreQueue.scala 164:59:@1860.6]
  assign _GEN_990 = _T_3637 ? 1'h1 : storeCompleted_15; // @[StoreQueue.scala 164:86:@1861.6]
  assign _GEN_991 = initBits_15 ? 1'h0 : _GEN_990; // @[StoreQueue.scala 162:37:@1854.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[StoreQueue.scala 180:72:@1865.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[StoreQueue.scala 180:72:@1867.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[StoreQueue.scala 180:72:@1869.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[StoreQueue.scala 180:72:@1871.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[StoreQueue.scala 180:72:@1873.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[StoreQueue.scala 180:72:@1875.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[StoreQueue.scala 180:72:@1877.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[StoreQueue.scala 180:72:@1879.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[StoreQueue.scala 180:72:@1881.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[StoreQueue.scala 180:72:@1883.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[StoreQueue.scala 180:72:@1885.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[StoreQueue.scala 180:72:@1887.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[StoreQueue.scala 180:72:@1889.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[StoreQueue.scala 180:72:@1891.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[StoreQueue.scala 180:72:@1893.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[StoreQueue.scala 180:72:@1895.4]
  assign _T_4122 = addrKnown_0 == 1'h0; // @[StoreQueue.scala 192:91:@1899.4]
  assign _T_4123 = entriesPorts_0_0 & _T_4122; // @[StoreQueue.scala 192:88:@1900.4]
  assign _T_4125 = addrKnown_1 == 1'h0; // @[StoreQueue.scala 192:91:@1901.4]
  assign _T_4126 = entriesPorts_0_1 & _T_4125; // @[StoreQueue.scala 192:88:@1902.4]
  assign _T_4128 = addrKnown_2 == 1'h0; // @[StoreQueue.scala 192:91:@1903.4]
  assign _T_4129 = entriesPorts_0_2 & _T_4128; // @[StoreQueue.scala 192:88:@1904.4]
  assign _T_4131 = addrKnown_3 == 1'h0; // @[StoreQueue.scala 192:91:@1905.4]
  assign _T_4132 = entriesPorts_0_3 & _T_4131; // @[StoreQueue.scala 192:88:@1906.4]
  assign _T_4134 = addrKnown_4 == 1'h0; // @[StoreQueue.scala 192:91:@1907.4]
  assign _T_4135 = entriesPorts_0_4 & _T_4134; // @[StoreQueue.scala 192:88:@1908.4]
  assign _T_4137 = addrKnown_5 == 1'h0; // @[StoreQueue.scala 192:91:@1909.4]
  assign _T_4138 = entriesPorts_0_5 & _T_4137; // @[StoreQueue.scala 192:88:@1910.4]
  assign _T_4140 = addrKnown_6 == 1'h0; // @[StoreQueue.scala 192:91:@1911.4]
  assign _T_4141 = entriesPorts_0_6 & _T_4140; // @[StoreQueue.scala 192:88:@1912.4]
  assign _T_4143 = addrKnown_7 == 1'h0; // @[StoreQueue.scala 192:91:@1913.4]
  assign _T_4144 = entriesPorts_0_7 & _T_4143; // @[StoreQueue.scala 192:88:@1914.4]
  assign _T_4146 = addrKnown_8 == 1'h0; // @[StoreQueue.scala 192:91:@1915.4]
  assign _T_4147 = entriesPorts_0_8 & _T_4146; // @[StoreQueue.scala 192:88:@1916.4]
  assign _T_4149 = addrKnown_9 == 1'h0; // @[StoreQueue.scala 192:91:@1917.4]
  assign _T_4150 = entriesPorts_0_9 & _T_4149; // @[StoreQueue.scala 192:88:@1918.4]
  assign _T_4152 = addrKnown_10 == 1'h0; // @[StoreQueue.scala 192:91:@1919.4]
  assign _T_4153 = entriesPorts_0_10 & _T_4152; // @[StoreQueue.scala 192:88:@1920.4]
  assign _T_4155 = addrKnown_11 == 1'h0; // @[StoreQueue.scala 192:91:@1921.4]
  assign _T_4156 = entriesPorts_0_11 & _T_4155; // @[StoreQueue.scala 192:88:@1922.4]
  assign _T_4158 = addrKnown_12 == 1'h0; // @[StoreQueue.scala 192:91:@1923.4]
  assign _T_4159 = entriesPorts_0_12 & _T_4158; // @[StoreQueue.scala 192:88:@1924.4]
  assign _T_4161 = addrKnown_13 == 1'h0; // @[StoreQueue.scala 192:91:@1925.4]
  assign _T_4162 = entriesPorts_0_13 & _T_4161; // @[StoreQueue.scala 192:88:@1926.4]
  assign _T_4164 = addrKnown_14 == 1'h0; // @[StoreQueue.scala 192:91:@1927.4]
  assign _T_4165 = entriesPorts_0_14 & _T_4164; // @[StoreQueue.scala 192:88:@1928.4]
  assign _T_4167 = addrKnown_15 == 1'h0; // @[StoreQueue.scala 192:91:@1929.4]
  assign _T_4168 = entriesPorts_0_15 & _T_4167; // @[StoreQueue.scala 192:88:@1930.4]
  assign _T_4192 = dataKnown_0 == 1'h0; // @[StoreQueue.scala 193:91:@1948.4]
  assign _T_4193 = entriesPorts_0_0 & _T_4192; // @[StoreQueue.scala 193:88:@1949.4]
  assign _T_4195 = dataKnown_1 == 1'h0; // @[StoreQueue.scala 193:91:@1950.4]
  assign _T_4196 = entriesPorts_0_1 & _T_4195; // @[StoreQueue.scala 193:88:@1951.4]
  assign _T_4198 = dataKnown_2 == 1'h0; // @[StoreQueue.scala 193:91:@1952.4]
  assign _T_4199 = entriesPorts_0_2 & _T_4198; // @[StoreQueue.scala 193:88:@1953.4]
  assign _T_4201 = dataKnown_3 == 1'h0; // @[StoreQueue.scala 193:91:@1954.4]
  assign _T_4202 = entriesPorts_0_3 & _T_4201; // @[StoreQueue.scala 193:88:@1955.4]
  assign _T_4204 = dataKnown_4 == 1'h0; // @[StoreQueue.scala 193:91:@1956.4]
  assign _T_4205 = entriesPorts_0_4 & _T_4204; // @[StoreQueue.scala 193:88:@1957.4]
  assign _T_4207 = dataKnown_5 == 1'h0; // @[StoreQueue.scala 193:91:@1958.4]
  assign _T_4208 = entriesPorts_0_5 & _T_4207; // @[StoreQueue.scala 193:88:@1959.4]
  assign _T_4210 = dataKnown_6 == 1'h0; // @[StoreQueue.scala 193:91:@1960.4]
  assign _T_4211 = entriesPorts_0_6 & _T_4210; // @[StoreQueue.scala 193:88:@1961.4]
  assign _T_4213 = dataKnown_7 == 1'h0; // @[StoreQueue.scala 193:91:@1962.4]
  assign _T_4214 = entriesPorts_0_7 & _T_4213; // @[StoreQueue.scala 193:88:@1963.4]
  assign _T_4216 = dataKnown_8 == 1'h0; // @[StoreQueue.scala 193:91:@1964.4]
  assign _T_4217 = entriesPorts_0_8 & _T_4216; // @[StoreQueue.scala 193:88:@1965.4]
  assign _T_4219 = dataKnown_9 == 1'h0; // @[StoreQueue.scala 193:91:@1966.4]
  assign _T_4220 = entriesPorts_0_9 & _T_4219; // @[StoreQueue.scala 193:88:@1967.4]
  assign _T_4222 = dataKnown_10 == 1'h0; // @[StoreQueue.scala 193:91:@1968.4]
  assign _T_4223 = entriesPorts_0_10 & _T_4222; // @[StoreQueue.scala 193:88:@1969.4]
  assign _T_4225 = dataKnown_11 == 1'h0; // @[StoreQueue.scala 193:91:@1970.4]
  assign _T_4226 = entriesPorts_0_11 & _T_4225; // @[StoreQueue.scala 193:88:@1971.4]
  assign _T_4228 = dataKnown_12 == 1'h0; // @[StoreQueue.scala 193:91:@1972.4]
  assign _T_4229 = entriesPorts_0_12 & _T_4228; // @[StoreQueue.scala 193:88:@1973.4]
  assign _T_4231 = dataKnown_13 == 1'h0; // @[StoreQueue.scala 193:91:@1974.4]
  assign _T_4232 = entriesPorts_0_13 & _T_4231; // @[StoreQueue.scala 193:88:@1975.4]
  assign _T_4234 = dataKnown_14 == 1'h0; // @[StoreQueue.scala 193:91:@1976.4]
  assign _T_4235 = entriesPorts_0_14 & _T_4234; // @[StoreQueue.scala 193:88:@1977.4]
  assign _T_4237 = dataKnown_15 == 1'h0; // @[StoreQueue.scala 193:91:@1978.4]
  assign _T_4238 = entriesPorts_0_15 & _T_4237; // @[StoreQueue.scala 193:88:@1979.4]
  assign _T_4263 = 16'h1 << head; // @[OneHot.scala 52:12:@1998.4]
  assign _T_4265 = _T_4263[0]; // @[util.scala 33:60:@2000.4]
  assign _T_4266 = _T_4263[1]; // @[util.scala 33:60:@2001.4]
  assign _T_4267 = _T_4263[2]; // @[util.scala 33:60:@2002.4]
  assign _T_4268 = _T_4263[3]; // @[util.scala 33:60:@2003.4]
  assign _T_4269 = _T_4263[4]; // @[util.scala 33:60:@2004.4]
  assign _T_4270 = _T_4263[5]; // @[util.scala 33:60:@2005.4]
  assign _T_4271 = _T_4263[6]; // @[util.scala 33:60:@2006.4]
  assign _T_4272 = _T_4263[7]; // @[util.scala 33:60:@2007.4]
  assign _T_4273 = _T_4263[8]; // @[util.scala 33:60:@2008.4]
  assign _T_4274 = _T_4263[9]; // @[util.scala 33:60:@2009.4]
  assign _T_4275 = _T_4263[10]; // @[util.scala 33:60:@2010.4]
  assign _T_4276 = _T_4263[11]; // @[util.scala 33:60:@2011.4]
  assign _T_4277 = _T_4263[12]; // @[util.scala 33:60:@2012.4]
  assign _T_4278 = _T_4263[13]; // @[util.scala 33:60:@2013.4]
  assign _T_4279 = _T_4263[14]; // @[util.scala 33:60:@2014.4]
  assign _T_4280 = _T_4263[15]; // @[util.scala 33:60:@2015.4]
  assign _T_4321 = _T_4168 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2033.4]
  assign _T_4322 = _T_4165 ? 16'h4000 : _T_4321; // @[Mux.scala 31:69:@2034.4]
  assign _T_4323 = _T_4162 ? 16'h2000 : _T_4322; // @[Mux.scala 31:69:@2035.4]
  assign _T_4324 = _T_4159 ? 16'h1000 : _T_4323; // @[Mux.scala 31:69:@2036.4]
  assign _T_4325 = _T_4156 ? 16'h800 : _T_4324; // @[Mux.scala 31:69:@2037.4]
  assign _T_4326 = _T_4153 ? 16'h400 : _T_4325; // @[Mux.scala 31:69:@2038.4]
  assign _T_4327 = _T_4150 ? 16'h200 : _T_4326; // @[Mux.scala 31:69:@2039.4]
  assign _T_4328 = _T_4147 ? 16'h100 : _T_4327; // @[Mux.scala 31:69:@2040.4]
  assign _T_4329 = _T_4144 ? 16'h80 : _T_4328; // @[Mux.scala 31:69:@2041.4]
  assign _T_4330 = _T_4141 ? 16'h40 : _T_4329; // @[Mux.scala 31:69:@2042.4]
  assign _T_4331 = _T_4138 ? 16'h20 : _T_4330; // @[Mux.scala 31:69:@2043.4]
  assign _T_4332 = _T_4135 ? 16'h10 : _T_4331; // @[Mux.scala 31:69:@2044.4]
  assign _T_4333 = _T_4132 ? 16'h8 : _T_4332; // @[Mux.scala 31:69:@2045.4]
  assign _T_4334 = _T_4129 ? 16'h4 : _T_4333; // @[Mux.scala 31:69:@2046.4]
  assign _T_4335 = _T_4126 ? 16'h2 : _T_4334; // @[Mux.scala 31:69:@2047.4]
  assign _T_4336 = _T_4123 ? 16'h1 : _T_4335; // @[Mux.scala 31:69:@2048.4]
  assign _T_4337 = _T_4336[0]; // @[OneHot.scala 66:30:@2049.4]
  assign _T_4338 = _T_4336[1]; // @[OneHot.scala 66:30:@2050.4]
  assign _T_4339 = _T_4336[2]; // @[OneHot.scala 66:30:@2051.4]
  assign _T_4340 = _T_4336[3]; // @[OneHot.scala 66:30:@2052.4]
  assign _T_4341 = _T_4336[4]; // @[OneHot.scala 66:30:@2053.4]
  assign _T_4342 = _T_4336[5]; // @[OneHot.scala 66:30:@2054.4]
  assign _T_4343 = _T_4336[6]; // @[OneHot.scala 66:30:@2055.4]
  assign _T_4344 = _T_4336[7]; // @[OneHot.scala 66:30:@2056.4]
  assign _T_4345 = _T_4336[8]; // @[OneHot.scala 66:30:@2057.4]
  assign _T_4346 = _T_4336[9]; // @[OneHot.scala 66:30:@2058.4]
  assign _T_4347 = _T_4336[10]; // @[OneHot.scala 66:30:@2059.4]
  assign _T_4348 = _T_4336[11]; // @[OneHot.scala 66:30:@2060.4]
  assign _T_4349 = _T_4336[12]; // @[OneHot.scala 66:30:@2061.4]
  assign _T_4350 = _T_4336[13]; // @[OneHot.scala 66:30:@2062.4]
  assign _T_4351 = _T_4336[14]; // @[OneHot.scala 66:30:@2063.4]
  assign _T_4352 = _T_4336[15]; // @[OneHot.scala 66:30:@2064.4]
  assign _T_4393 = _T_4123 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2082.4]
  assign _T_4394 = _T_4168 ? 16'h4000 : _T_4393; // @[Mux.scala 31:69:@2083.4]
  assign _T_4395 = _T_4165 ? 16'h2000 : _T_4394; // @[Mux.scala 31:69:@2084.4]
  assign _T_4396 = _T_4162 ? 16'h1000 : _T_4395; // @[Mux.scala 31:69:@2085.4]
  assign _T_4397 = _T_4159 ? 16'h800 : _T_4396; // @[Mux.scala 31:69:@2086.4]
  assign _T_4398 = _T_4156 ? 16'h400 : _T_4397; // @[Mux.scala 31:69:@2087.4]
  assign _T_4399 = _T_4153 ? 16'h200 : _T_4398; // @[Mux.scala 31:69:@2088.4]
  assign _T_4400 = _T_4150 ? 16'h100 : _T_4399; // @[Mux.scala 31:69:@2089.4]
  assign _T_4401 = _T_4147 ? 16'h80 : _T_4400; // @[Mux.scala 31:69:@2090.4]
  assign _T_4402 = _T_4144 ? 16'h40 : _T_4401; // @[Mux.scala 31:69:@2091.4]
  assign _T_4403 = _T_4141 ? 16'h20 : _T_4402; // @[Mux.scala 31:69:@2092.4]
  assign _T_4404 = _T_4138 ? 16'h10 : _T_4403; // @[Mux.scala 31:69:@2093.4]
  assign _T_4405 = _T_4135 ? 16'h8 : _T_4404; // @[Mux.scala 31:69:@2094.4]
  assign _T_4406 = _T_4132 ? 16'h4 : _T_4405; // @[Mux.scala 31:69:@2095.4]
  assign _T_4407 = _T_4129 ? 16'h2 : _T_4406; // @[Mux.scala 31:69:@2096.4]
  assign _T_4408 = _T_4126 ? 16'h1 : _T_4407; // @[Mux.scala 31:69:@2097.4]
  assign _T_4409 = _T_4408[0]; // @[OneHot.scala 66:30:@2098.4]
  assign _T_4410 = _T_4408[1]; // @[OneHot.scala 66:30:@2099.4]
  assign _T_4411 = _T_4408[2]; // @[OneHot.scala 66:30:@2100.4]
  assign _T_4412 = _T_4408[3]; // @[OneHot.scala 66:30:@2101.4]
  assign _T_4413 = _T_4408[4]; // @[OneHot.scala 66:30:@2102.4]
  assign _T_4414 = _T_4408[5]; // @[OneHot.scala 66:30:@2103.4]
  assign _T_4415 = _T_4408[6]; // @[OneHot.scala 66:30:@2104.4]
  assign _T_4416 = _T_4408[7]; // @[OneHot.scala 66:30:@2105.4]
  assign _T_4417 = _T_4408[8]; // @[OneHot.scala 66:30:@2106.4]
  assign _T_4418 = _T_4408[9]; // @[OneHot.scala 66:30:@2107.4]
  assign _T_4419 = _T_4408[10]; // @[OneHot.scala 66:30:@2108.4]
  assign _T_4420 = _T_4408[11]; // @[OneHot.scala 66:30:@2109.4]
  assign _T_4421 = _T_4408[12]; // @[OneHot.scala 66:30:@2110.4]
  assign _T_4422 = _T_4408[13]; // @[OneHot.scala 66:30:@2111.4]
  assign _T_4423 = _T_4408[14]; // @[OneHot.scala 66:30:@2112.4]
  assign _T_4424 = _T_4408[15]; // @[OneHot.scala 66:30:@2113.4]
  assign _T_4465 = _T_4126 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2131.4]
  assign _T_4466 = _T_4123 ? 16'h4000 : _T_4465; // @[Mux.scala 31:69:@2132.4]
  assign _T_4467 = _T_4168 ? 16'h2000 : _T_4466; // @[Mux.scala 31:69:@2133.4]
  assign _T_4468 = _T_4165 ? 16'h1000 : _T_4467; // @[Mux.scala 31:69:@2134.4]
  assign _T_4469 = _T_4162 ? 16'h800 : _T_4468; // @[Mux.scala 31:69:@2135.4]
  assign _T_4470 = _T_4159 ? 16'h400 : _T_4469; // @[Mux.scala 31:69:@2136.4]
  assign _T_4471 = _T_4156 ? 16'h200 : _T_4470; // @[Mux.scala 31:69:@2137.4]
  assign _T_4472 = _T_4153 ? 16'h100 : _T_4471; // @[Mux.scala 31:69:@2138.4]
  assign _T_4473 = _T_4150 ? 16'h80 : _T_4472; // @[Mux.scala 31:69:@2139.4]
  assign _T_4474 = _T_4147 ? 16'h40 : _T_4473; // @[Mux.scala 31:69:@2140.4]
  assign _T_4475 = _T_4144 ? 16'h20 : _T_4474; // @[Mux.scala 31:69:@2141.4]
  assign _T_4476 = _T_4141 ? 16'h10 : _T_4475; // @[Mux.scala 31:69:@2142.4]
  assign _T_4477 = _T_4138 ? 16'h8 : _T_4476; // @[Mux.scala 31:69:@2143.4]
  assign _T_4478 = _T_4135 ? 16'h4 : _T_4477; // @[Mux.scala 31:69:@2144.4]
  assign _T_4479 = _T_4132 ? 16'h2 : _T_4478; // @[Mux.scala 31:69:@2145.4]
  assign _T_4480 = _T_4129 ? 16'h1 : _T_4479; // @[Mux.scala 31:69:@2146.4]
  assign _T_4481 = _T_4480[0]; // @[OneHot.scala 66:30:@2147.4]
  assign _T_4482 = _T_4480[1]; // @[OneHot.scala 66:30:@2148.4]
  assign _T_4483 = _T_4480[2]; // @[OneHot.scala 66:30:@2149.4]
  assign _T_4484 = _T_4480[3]; // @[OneHot.scala 66:30:@2150.4]
  assign _T_4485 = _T_4480[4]; // @[OneHot.scala 66:30:@2151.4]
  assign _T_4486 = _T_4480[5]; // @[OneHot.scala 66:30:@2152.4]
  assign _T_4487 = _T_4480[6]; // @[OneHot.scala 66:30:@2153.4]
  assign _T_4488 = _T_4480[7]; // @[OneHot.scala 66:30:@2154.4]
  assign _T_4489 = _T_4480[8]; // @[OneHot.scala 66:30:@2155.4]
  assign _T_4490 = _T_4480[9]; // @[OneHot.scala 66:30:@2156.4]
  assign _T_4491 = _T_4480[10]; // @[OneHot.scala 66:30:@2157.4]
  assign _T_4492 = _T_4480[11]; // @[OneHot.scala 66:30:@2158.4]
  assign _T_4493 = _T_4480[12]; // @[OneHot.scala 66:30:@2159.4]
  assign _T_4494 = _T_4480[13]; // @[OneHot.scala 66:30:@2160.4]
  assign _T_4495 = _T_4480[14]; // @[OneHot.scala 66:30:@2161.4]
  assign _T_4496 = _T_4480[15]; // @[OneHot.scala 66:30:@2162.4]
  assign _T_4537 = _T_4129 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2180.4]
  assign _T_4538 = _T_4126 ? 16'h4000 : _T_4537; // @[Mux.scala 31:69:@2181.4]
  assign _T_4539 = _T_4123 ? 16'h2000 : _T_4538; // @[Mux.scala 31:69:@2182.4]
  assign _T_4540 = _T_4168 ? 16'h1000 : _T_4539; // @[Mux.scala 31:69:@2183.4]
  assign _T_4541 = _T_4165 ? 16'h800 : _T_4540; // @[Mux.scala 31:69:@2184.4]
  assign _T_4542 = _T_4162 ? 16'h400 : _T_4541; // @[Mux.scala 31:69:@2185.4]
  assign _T_4543 = _T_4159 ? 16'h200 : _T_4542; // @[Mux.scala 31:69:@2186.4]
  assign _T_4544 = _T_4156 ? 16'h100 : _T_4543; // @[Mux.scala 31:69:@2187.4]
  assign _T_4545 = _T_4153 ? 16'h80 : _T_4544; // @[Mux.scala 31:69:@2188.4]
  assign _T_4546 = _T_4150 ? 16'h40 : _T_4545; // @[Mux.scala 31:69:@2189.4]
  assign _T_4547 = _T_4147 ? 16'h20 : _T_4546; // @[Mux.scala 31:69:@2190.4]
  assign _T_4548 = _T_4144 ? 16'h10 : _T_4547; // @[Mux.scala 31:69:@2191.4]
  assign _T_4549 = _T_4141 ? 16'h8 : _T_4548; // @[Mux.scala 31:69:@2192.4]
  assign _T_4550 = _T_4138 ? 16'h4 : _T_4549; // @[Mux.scala 31:69:@2193.4]
  assign _T_4551 = _T_4135 ? 16'h2 : _T_4550; // @[Mux.scala 31:69:@2194.4]
  assign _T_4552 = _T_4132 ? 16'h1 : _T_4551; // @[Mux.scala 31:69:@2195.4]
  assign _T_4553 = _T_4552[0]; // @[OneHot.scala 66:30:@2196.4]
  assign _T_4554 = _T_4552[1]; // @[OneHot.scala 66:30:@2197.4]
  assign _T_4555 = _T_4552[2]; // @[OneHot.scala 66:30:@2198.4]
  assign _T_4556 = _T_4552[3]; // @[OneHot.scala 66:30:@2199.4]
  assign _T_4557 = _T_4552[4]; // @[OneHot.scala 66:30:@2200.4]
  assign _T_4558 = _T_4552[5]; // @[OneHot.scala 66:30:@2201.4]
  assign _T_4559 = _T_4552[6]; // @[OneHot.scala 66:30:@2202.4]
  assign _T_4560 = _T_4552[7]; // @[OneHot.scala 66:30:@2203.4]
  assign _T_4561 = _T_4552[8]; // @[OneHot.scala 66:30:@2204.4]
  assign _T_4562 = _T_4552[9]; // @[OneHot.scala 66:30:@2205.4]
  assign _T_4563 = _T_4552[10]; // @[OneHot.scala 66:30:@2206.4]
  assign _T_4564 = _T_4552[11]; // @[OneHot.scala 66:30:@2207.4]
  assign _T_4565 = _T_4552[12]; // @[OneHot.scala 66:30:@2208.4]
  assign _T_4566 = _T_4552[13]; // @[OneHot.scala 66:30:@2209.4]
  assign _T_4567 = _T_4552[14]; // @[OneHot.scala 66:30:@2210.4]
  assign _T_4568 = _T_4552[15]; // @[OneHot.scala 66:30:@2211.4]
  assign _T_4609 = _T_4132 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2229.4]
  assign _T_4610 = _T_4129 ? 16'h4000 : _T_4609; // @[Mux.scala 31:69:@2230.4]
  assign _T_4611 = _T_4126 ? 16'h2000 : _T_4610; // @[Mux.scala 31:69:@2231.4]
  assign _T_4612 = _T_4123 ? 16'h1000 : _T_4611; // @[Mux.scala 31:69:@2232.4]
  assign _T_4613 = _T_4168 ? 16'h800 : _T_4612; // @[Mux.scala 31:69:@2233.4]
  assign _T_4614 = _T_4165 ? 16'h400 : _T_4613; // @[Mux.scala 31:69:@2234.4]
  assign _T_4615 = _T_4162 ? 16'h200 : _T_4614; // @[Mux.scala 31:69:@2235.4]
  assign _T_4616 = _T_4159 ? 16'h100 : _T_4615; // @[Mux.scala 31:69:@2236.4]
  assign _T_4617 = _T_4156 ? 16'h80 : _T_4616; // @[Mux.scala 31:69:@2237.4]
  assign _T_4618 = _T_4153 ? 16'h40 : _T_4617; // @[Mux.scala 31:69:@2238.4]
  assign _T_4619 = _T_4150 ? 16'h20 : _T_4618; // @[Mux.scala 31:69:@2239.4]
  assign _T_4620 = _T_4147 ? 16'h10 : _T_4619; // @[Mux.scala 31:69:@2240.4]
  assign _T_4621 = _T_4144 ? 16'h8 : _T_4620; // @[Mux.scala 31:69:@2241.4]
  assign _T_4622 = _T_4141 ? 16'h4 : _T_4621; // @[Mux.scala 31:69:@2242.4]
  assign _T_4623 = _T_4138 ? 16'h2 : _T_4622; // @[Mux.scala 31:69:@2243.4]
  assign _T_4624 = _T_4135 ? 16'h1 : _T_4623; // @[Mux.scala 31:69:@2244.4]
  assign _T_4625 = _T_4624[0]; // @[OneHot.scala 66:30:@2245.4]
  assign _T_4626 = _T_4624[1]; // @[OneHot.scala 66:30:@2246.4]
  assign _T_4627 = _T_4624[2]; // @[OneHot.scala 66:30:@2247.4]
  assign _T_4628 = _T_4624[3]; // @[OneHot.scala 66:30:@2248.4]
  assign _T_4629 = _T_4624[4]; // @[OneHot.scala 66:30:@2249.4]
  assign _T_4630 = _T_4624[5]; // @[OneHot.scala 66:30:@2250.4]
  assign _T_4631 = _T_4624[6]; // @[OneHot.scala 66:30:@2251.4]
  assign _T_4632 = _T_4624[7]; // @[OneHot.scala 66:30:@2252.4]
  assign _T_4633 = _T_4624[8]; // @[OneHot.scala 66:30:@2253.4]
  assign _T_4634 = _T_4624[9]; // @[OneHot.scala 66:30:@2254.4]
  assign _T_4635 = _T_4624[10]; // @[OneHot.scala 66:30:@2255.4]
  assign _T_4636 = _T_4624[11]; // @[OneHot.scala 66:30:@2256.4]
  assign _T_4637 = _T_4624[12]; // @[OneHot.scala 66:30:@2257.4]
  assign _T_4638 = _T_4624[13]; // @[OneHot.scala 66:30:@2258.4]
  assign _T_4639 = _T_4624[14]; // @[OneHot.scala 66:30:@2259.4]
  assign _T_4640 = _T_4624[15]; // @[OneHot.scala 66:30:@2260.4]
  assign _T_4681 = _T_4135 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2278.4]
  assign _T_4682 = _T_4132 ? 16'h4000 : _T_4681; // @[Mux.scala 31:69:@2279.4]
  assign _T_4683 = _T_4129 ? 16'h2000 : _T_4682; // @[Mux.scala 31:69:@2280.4]
  assign _T_4684 = _T_4126 ? 16'h1000 : _T_4683; // @[Mux.scala 31:69:@2281.4]
  assign _T_4685 = _T_4123 ? 16'h800 : _T_4684; // @[Mux.scala 31:69:@2282.4]
  assign _T_4686 = _T_4168 ? 16'h400 : _T_4685; // @[Mux.scala 31:69:@2283.4]
  assign _T_4687 = _T_4165 ? 16'h200 : _T_4686; // @[Mux.scala 31:69:@2284.4]
  assign _T_4688 = _T_4162 ? 16'h100 : _T_4687; // @[Mux.scala 31:69:@2285.4]
  assign _T_4689 = _T_4159 ? 16'h80 : _T_4688; // @[Mux.scala 31:69:@2286.4]
  assign _T_4690 = _T_4156 ? 16'h40 : _T_4689; // @[Mux.scala 31:69:@2287.4]
  assign _T_4691 = _T_4153 ? 16'h20 : _T_4690; // @[Mux.scala 31:69:@2288.4]
  assign _T_4692 = _T_4150 ? 16'h10 : _T_4691; // @[Mux.scala 31:69:@2289.4]
  assign _T_4693 = _T_4147 ? 16'h8 : _T_4692; // @[Mux.scala 31:69:@2290.4]
  assign _T_4694 = _T_4144 ? 16'h4 : _T_4693; // @[Mux.scala 31:69:@2291.4]
  assign _T_4695 = _T_4141 ? 16'h2 : _T_4694; // @[Mux.scala 31:69:@2292.4]
  assign _T_4696 = _T_4138 ? 16'h1 : _T_4695; // @[Mux.scala 31:69:@2293.4]
  assign _T_4697 = _T_4696[0]; // @[OneHot.scala 66:30:@2294.4]
  assign _T_4698 = _T_4696[1]; // @[OneHot.scala 66:30:@2295.4]
  assign _T_4699 = _T_4696[2]; // @[OneHot.scala 66:30:@2296.4]
  assign _T_4700 = _T_4696[3]; // @[OneHot.scala 66:30:@2297.4]
  assign _T_4701 = _T_4696[4]; // @[OneHot.scala 66:30:@2298.4]
  assign _T_4702 = _T_4696[5]; // @[OneHot.scala 66:30:@2299.4]
  assign _T_4703 = _T_4696[6]; // @[OneHot.scala 66:30:@2300.4]
  assign _T_4704 = _T_4696[7]; // @[OneHot.scala 66:30:@2301.4]
  assign _T_4705 = _T_4696[8]; // @[OneHot.scala 66:30:@2302.4]
  assign _T_4706 = _T_4696[9]; // @[OneHot.scala 66:30:@2303.4]
  assign _T_4707 = _T_4696[10]; // @[OneHot.scala 66:30:@2304.4]
  assign _T_4708 = _T_4696[11]; // @[OneHot.scala 66:30:@2305.4]
  assign _T_4709 = _T_4696[12]; // @[OneHot.scala 66:30:@2306.4]
  assign _T_4710 = _T_4696[13]; // @[OneHot.scala 66:30:@2307.4]
  assign _T_4711 = _T_4696[14]; // @[OneHot.scala 66:30:@2308.4]
  assign _T_4712 = _T_4696[15]; // @[OneHot.scala 66:30:@2309.4]
  assign _T_4753 = _T_4138 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2327.4]
  assign _T_4754 = _T_4135 ? 16'h4000 : _T_4753; // @[Mux.scala 31:69:@2328.4]
  assign _T_4755 = _T_4132 ? 16'h2000 : _T_4754; // @[Mux.scala 31:69:@2329.4]
  assign _T_4756 = _T_4129 ? 16'h1000 : _T_4755; // @[Mux.scala 31:69:@2330.4]
  assign _T_4757 = _T_4126 ? 16'h800 : _T_4756; // @[Mux.scala 31:69:@2331.4]
  assign _T_4758 = _T_4123 ? 16'h400 : _T_4757; // @[Mux.scala 31:69:@2332.4]
  assign _T_4759 = _T_4168 ? 16'h200 : _T_4758; // @[Mux.scala 31:69:@2333.4]
  assign _T_4760 = _T_4165 ? 16'h100 : _T_4759; // @[Mux.scala 31:69:@2334.4]
  assign _T_4761 = _T_4162 ? 16'h80 : _T_4760; // @[Mux.scala 31:69:@2335.4]
  assign _T_4762 = _T_4159 ? 16'h40 : _T_4761; // @[Mux.scala 31:69:@2336.4]
  assign _T_4763 = _T_4156 ? 16'h20 : _T_4762; // @[Mux.scala 31:69:@2337.4]
  assign _T_4764 = _T_4153 ? 16'h10 : _T_4763; // @[Mux.scala 31:69:@2338.4]
  assign _T_4765 = _T_4150 ? 16'h8 : _T_4764; // @[Mux.scala 31:69:@2339.4]
  assign _T_4766 = _T_4147 ? 16'h4 : _T_4765; // @[Mux.scala 31:69:@2340.4]
  assign _T_4767 = _T_4144 ? 16'h2 : _T_4766; // @[Mux.scala 31:69:@2341.4]
  assign _T_4768 = _T_4141 ? 16'h1 : _T_4767; // @[Mux.scala 31:69:@2342.4]
  assign _T_4769 = _T_4768[0]; // @[OneHot.scala 66:30:@2343.4]
  assign _T_4770 = _T_4768[1]; // @[OneHot.scala 66:30:@2344.4]
  assign _T_4771 = _T_4768[2]; // @[OneHot.scala 66:30:@2345.4]
  assign _T_4772 = _T_4768[3]; // @[OneHot.scala 66:30:@2346.4]
  assign _T_4773 = _T_4768[4]; // @[OneHot.scala 66:30:@2347.4]
  assign _T_4774 = _T_4768[5]; // @[OneHot.scala 66:30:@2348.4]
  assign _T_4775 = _T_4768[6]; // @[OneHot.scala 66:30:@2349.4]
  assign _T_4776 = _T_4768[7]; // @[OneHot.scala 66:30:@2350.4]
  assign _T_4777 = _T_4768[8]; // @[OneHot.scala 66:30:@2351.4]
  assign _T_4778 = _T_4768[9]; // @[OneHot.scala 66:30:@2352.4]
  assign _T_4779 = _T_4768[10]; // @[OneHot.scala 66:30:@2353.4]
  assign _T_4780 = _T_4768[11]; // @[OneHot.scala 66:30:@2354.4]
  assign _T_4781 = _T_4768[12]; // @[OneHot.scala 66:30:@2355.4]
  assign _T_4782 = _T_4768[13]; // @[OneHot.scala 66:30:@2356.4]
  assign _T_4783 = _T_4768[14]; // @[OneHot.scala 66:30:@2357.4]
  assign _T_4784 = _T_4768[15]; // @[OneHot.scala 66:30:@2358.4]
  assign _T_4825 = _T_4141 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2376.4]
  assign _T_4826 = _T_4138 ? 16'h4000 : _T_4825; // @[Mux.scala 31:69:@2377.4]
  assign _T_4827 = _T_4135 ? 16'h2000 : _T_4826; // @[Mux.scala 31:69:@2378.4]
  assign _T_4828 = _T_4132 ? 16'h1000 : _T_4827; // @[Mux.scala 31:69:@2379.4]
  assign _T_4829 = _T_4129 ? 16'h800 : _T_4828; // @[Mux.scala 31:69:@2380.4]
  assign _T_4830 = _T_4126 ? 16'h400 : _T_4829; // @[Mux.scala 31:69:@2381.4]
  assign _T_4831 = _T_4123 ? 16'h200 : _T_4830; // @[Mux.scala 31:69:@2382.4]
  assign _T_4832 = _T_4168 ? 16'h100 : _T_4831; // @[Mux.scala 31:69:@2383.4]
  assign _T_4833 = _T_4165 ? 16'h80 : _T_4832; // @[Mux.scala 31:69:@2384.4]
  assign _T_4834 = _T_4162 ? 16'h40 : _T_4833; // @[Mux.scala 31:69:@2385.4]
  assign _T_4835 = _T_4159 ? 16'h20 : _T_4834; // @[Mux.scala 31:69:@2386.4]
  assign _T_4836 = _T_4156 ? 16'h10 : _T_4835; // @[Mux.scala 31:69:@2387.4]
  assign _T_4837 = _T_4153 ? 16'h8 : _T_4836; // @[Mux.scala 31:69:@2388.4]
  assign _T_4838 = _T_4150 ? 16'h4 : _T_4837; // @[Mux.scala 31:69:@2389.4]
  assign _T_4839 = _T_4147 ? 16'h2 : _T_4838; // @[Mux.scala 31:69:@2390.4]
  assign _T_4840 = _T_4144 ? 16'h1 : _T_4839; // @[Mux.scala 31:69:@2391.4]
  assign _T_4841 = _T_4840[0]; // @[OneHot.scala 66:30:@2392.4]
  assign _T_4842 = _T_4840[1]; // @[OneHot.scala 66:30:@2393.4]
  assign _T_4843 = _T_4840[2]; // @[OneHot.scala 66:30:@2394.4]
  assign _T_4844 = _T_4840[3]; // @[OneHot.scala 66:30:@2395.4]
  assign _T_4845 = _T_4840[4]; // @[OneHot.scala 66:30:@2396.4]
  assign _T_4846 = _T_4840[5]; // @[OneHot.scala 66:30:@2397.4]
  assign _T_4847 = _T_4840[6]; // @[OneHot.scala 66:30:@2398.4]
  assign _T_4848 = _T_4840[7]; // @[OneHot.scala 66:30:@2399.4]
  assign _T_4849 = _T_4840[8]; // @[OneHot.scala 66:30:@2400.4]
  assign _T_4850 = _T_4840[9]; // @[OneHot.scala 66:30:@2401.4]
  assign _T_4851 = _T_4840[10]; // @[OneHot.scala 66:30:@2402.4]
  assign _T_4852 = _T_4840[11]; // @[OneHot.scala 66:30:@2403.4]
  assign _T_4853 = _T_4840[12]; // @[OneHot.scala 66:30:@2404.4]
  assign _T_4854 = _T_4840[13]; // @[OneHot.scala 66:30:@2405.4]
  assign _T_4855 = _T_4840[14]; // @[OneHot.scala 66:30:@2406.4]
  assign _T_4856 = _T_4840[15]; // @[OneHot.scala 66:30:@2407.4]
  assign _T_4897 = _T_4144 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2425.4]
  assign _T_4898 = _T_4141 ? 16'h4000 : _T_4897; // @[Mux.scala 31:69:@2426.4]
  assign _T_4899 = _T_4138 ? 16'h2000 : _T_4898; // @[Mux.scala 31:69:@2427.4]
  assign _T_4900 = _T_4135 ? 16'h1000 : _T_4899; // @[Mux.scala 31:69:@2428.4]
  assign _T_4901 = _T_4132 ? 16'h800 : _T_4900; // @[Mux.scala 31:69:@2429.4]
  assign _T_4902 = _T_4129 ? 16'h400 : _T_4901; // @[Mux.scala 31:69:@2430.4]
  assign _T_4903 = _T_4126 ? 16'h200 : _T_4902; // @[Mux.scala 31:69:@2431.4]
  assign _T_4904 = _T_4123 ? 16'h100 : _T_4903; // @[Mux.scala 31:69:@2432.4]
  assign _T_4905 = _T_4168 ? 16'h80 : _T_4904; // @[Mux.scala 31:69:@2433.4]
  assign _T_4906 = _T_4165 ? 16'h40 : _T_4905; // @[Mux.scala 31:69:@2434.4]
  assign _T_4907 = _T_4162 ? 16'h20 : _T_4906; // @[Mux.scala 31:69:@2435.4]
  assign _T_4908 = _T_4159 ? 16'h10 : _T_4907; // @[Mux.scala 31:69:@2436.4]
  assign _T_4909 = _T_4156 ? 16'h8 : _T_4908; // @[Mux.scala 31:69:@2437.4]
  assign _T_4910 = _T_4153 ? 16'h4 : _T_4909; // @[Mux.scala 31:69:@2438.4]
  assign _T_4911 = _T_4150 ? 16'h2 : _T_4910; // @[Mux.scala 31:69:@2439.4]
  assign _T_4912 = _T_4147 ? 16'h1 : _T_4911; // @[Mux.scala 31:69:@2440.4]
  assign _T_4913 = _T_4912[0]; // @[OneHot.scala 66:30:@2441.4]
  assign _T_4914 = _T_4912[1]; // @[OneHot.scala 66:30:@2442.4]
  assign _T_4915 = _T_4912[2]; // @[OneHot.scala 66:30:@2443.4]
  assign _T_4916 = _T_4912[3]; // @[OneHot.scala 66:30:@2444.4]
  assign _T_4917 = _T_4912[4]; // @[OneHot.scala 66:30:@2445.4]
  assign _T_4918 = _T_4912[5]; // @[OneHot.scala 66:30:@2446.4]
  assign _T_4919 = _T_4912[6]; // @[OneHot.scala 66:30:@2447.4]
  assign _T_4920 = _T_4912[7]; // @[OneHot.scala 66:30:@2448.4]
  assign _T_4921 = _T_4912[8]; // @[OneHot.scala 66:30:@2449.4]
  assign _T_4922 = _T_4912[9]; // @[OneHot.scala 66:30:@2450.4]
  assign _T_4923 = _T_4912[10]; // @[OneHot.scala 66:30:@2451.4]
  assign _T_4924 = _T_4912[11]; // @[OneHot.scala 66:30:@2452.4]
  assign _T_4925 = _T_4912[12]; // @[OneHot.scala 66:30:@2453.4]
  assign _T_4926 = _T_4912[13]; // @[OneHot.scala 66:30:@2454.4]
  assign _T_4927 = _T_4912[14]; // @[OneHot.scala 66:30:@2455.4]
  assign _T_4928 = _T_4912[15]; // @[OneHot.scala 66:30:@2456.4]
  assign _T_4969 = _T_4147 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2474.4]
  assign _T_4970 = _T_4144 ? 16'h4000 : _T_4969; // @[Mux.scala 31:69:@2475.4]
  assign _T_4971 = _T_4141 ? 16'h2000 : _T_4970; // @[Mux.scala 31:69:@2476.4]
  assign _T_4972 = _T_4138 ? 16'h1000 : _T_4971; // @[Mux.scala 31:69:@2477.4]
  assign _T_4973 = _T_4135 ? 16'h800 : _T_4972; // @[Mux.scala 31:69:@2478.4]
  assign _T_4974 = _T_4132 ? 16'h400 : _T_4973; // @[Mux.scala 31:69:@2479.4]
  assign _T_4975 = _T_4129 ? 16'h200 : _T_4974; // @[Mux.scala 31:69:@2480.4]
  assign _T_4976 = _T_4126 ? 16'h100 : _T_4975; // @[Mux.scala 31:69:@2481.4]
  assign _T_4977 = _T_4123 ? 16'h80 : _T_4976; // @[Mux.scala 31:69:@2482.4]
  assign _T_4978 = _T_4168 ? 16'h40 : _T_4977; // @[Mux.scala 31:69:@2483.4]
  assign _T_4979 = _T_4165 ? 16'h20 : _T_4978; // @[Mux.scala 31:69:@2484.4]
  assign _T_4980 = _T_4162 ? 16'h10 : _T_4979; // @[Mux.scala 31:69:@2485.4]
  assign _T_4981 = _T_4159 ? 16'h8 : _T_4980; // @[Mux.scala 31:69:@2486.4]
  assign _T_4982 = _T_4156 ? 16'h4 : _T_4981; // @[Mux.scala 31:69:@2487.4]
  assign _T_4983 = _T_4153 ? 16'h2 : _T_4982; // @[Mux.scala 31:69:@2488.4]
  assign _T_4984 = _T_4150 ? 16'h1 : _T_4983; // @[Mux.scala 31:69:@2489.4]
  assign _T_4985 = _T_4984[0]; // @[OneHot.scala 66:30:@2490.4]
  assign _T_4986 = _T_4984[1]; // @[OneHot.scala 66:30:@2491.4]
  assign _T_4987 = _T_4984[2]; // @[OneHot.scala 66:30:@2492.4]
  assign _T_4988 = _T_4984[3]; // @[OneHot.scala 66:30:@2493.4]
  assign _T_4989 = _T_4984[4]; // @[OneHot.scala 66:30:@2494.4]
  assign _T_4990 = _T_4984[5]; // @[OneHot.scala 66:30:@2495.4]
  assign _T_4991 = _T_4984[6]; // @[OneHot.scala 66:30:@2496.4]
  assign _T_4992 = _T_4984[7]; // @[OneHot.scala 66:30:@2497.4]
  assign _T_4993 = _T_4984[8]; // @[OneHot.scala 66:30:@2498.4]
  assign _T_4994 = _T_4984[9]; // @[OneHot.scala 66:30:@2499.4]
  assign _T_4995 = _T_4984[10]; // @[OneHot.scala 66:30:@2500.4]
  assign _T_4996 = _T_4984[11]; // @[OneHot.scala 66:30:@2501.4]
  assign _T_4997 = _T_4984[12]; // @[OneHot.scala 66:30:@2502.4]
  assign _T_4998 = _T_4984[13]; // @[OneHot.scala 66:30:@2503.4]
  assign _T_4999 = _T_4984[14]; // @[OneHot.scala 66:30:@2504.4]
  assign _T_5000 = _T_4984[15]; // @[OneHot.scala 66:30:@2505.4]
  assign _T_5041 = _T_4150 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2523.4]
  assign _T_5042 = _T_4147 ? 16'h4000 : _T_5041; // @[Mux.scala 31:69:@2524.4]
  assign _T_5043 = _T_4144 ? 16'h2000 : _T_5042; // @[Mux.scala 31:69:@2525.4]
  assign _T_5044 = _T_4141 ? 16'h1000 : _T_5043; // @[Mux.scala 31:69:@2526.4]
  assign _T_5045 = _T_4138 ? 16'h800 : _T_5044; // @[Mux.scala 31:69:@2527.4]
  assign _T_5046 = _T_4135 ? 16'h400 : _T_5045; // @[Mux.scala 31:69:@2528.4]
  assign _T_5047 = _T_4132 ? 16'h200 : _T_5046; // @[Mux.scala 31:69:@2529.4]
  assign _T_5048 = _T_4129 ? 16'h100 : _T_5047; // @[Mux.scala 31:69:@2530.4]
  assign _T_5049 = _T_4126 ? 16'h80 : _T_5048; // @[Mux.scala 31:69:@2531.4]
  assign _T_5050 = _T_4123 ? 16'h40 : _T_5049; // @[Mux.scala 31:69:@2532.4]
  assign _T_5051 = _T_4168 ? 16'h20 : _T_5050; // @[Mux.scala 31:69:@2533.4]
  assign _T_5052 = _T_4165 ? 16'h10 : _T_5051; // @[Mux.scala 31:69:@2534.4]
  assign _T_5053 = _T_4162 ? 16'h8 : _T_5052; // @[Mux.scala 31:69:@2535.4]
  assign _T_5054 = _T_4159 ? 16'h4 : _T_5053; // @[Mux.scala 31:69:@2536.4]
  assign _T_5055 = _T_4156 ? 16'h2 : _T_5054; // @[Mux.scala 31:69:@2537.4]
  assign _T_5056 = _T_4153 ? 16'h1 : _T_5055; // @[Mux.scala 31:69:@2538.4]
  assign _T_5057 = _T_5056[0]; // @[OneHot.scala 66:30:@2539.4]
  assign _T_5058 = _T_5056[1]; // @[OneHot.scala 66:30:@2540.4]
  assign _T_5059 = _T_5056[2]; // @[OneHot.scala 66:30:@2541.4]
  assign _T_5060 = _T_5056[3]; // @[OneHot.scala 66:30:@2542.4]
  assign _T_5061 = _T_5056[4]; // @[OneHot.scala 66:30:@2543.4]
  assign _T_5062 = _T_5056[5]; // @[OneHot.scala 66:30:@2544.4]
  assign _T_5063 = _T_5056[6]; // @[OneHot.scala 66:30:@2545.4]
  assign _T_5064 = _T_5056[7]; // @[OneHot.scala 66:30:@2546.4]
  assign _T_5065 = _T_5056[8]; // @[OneHot.scala 66:30:@2547.4]
  assign _T_5066 = _T_5056[9]; // @[OneHot.scala 66:30:@2548.4]
  assign _T_5067 = _T_5056[10]; // @[OneHot.scala 66:30:@2549.4]
  assign _T_5068 = _T_5056[11]; // @[OneHot.scala 66:30:@2550.4]
  assign _T_5069 = _T_5056[12]; // @[OneHot.scala 66:30:@2551.4]
  assign _T_5070 = _T_5056[13]; // @[OneHot.scala 66:30:@2552.4]
  assign _T_5071 = _T_5056[14]; // @[OneHot.scala 66:30:@2553.4]
  assign _T_5072 = _T_5056[15]; // @[OneHot.scala 66:30:@2554.4]
  assign _T_5113 = _T_4153 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2572.4]
  assign _T_5114 = _T_4150 ? 16'h4000 : _T_5113; // @[Mux.scala 31:69:@2573.4]
  assign _T_5115 = _T_4147 ? 16'h2000 : _T_5114; // @[Mux.scala 31:69:@2574.4]
  assign _T_5116 = _T_4144 ? 16'h1000 : _T_5115; // @[Mux.scala 31:69:@2575.4]
  assign _T_5117 = _T_4141 ? 16'h800 : _T_5116; // @[Mux.scala 31:69:@2576.4]
  assign _T_5118 = _T_4138 ? 16'h400 : _T_5117; // @[Mux.scala 31:69:@2577.4]
  assign _T_5119 = _T_4135 ? 16'h200 : _T_5118; // @[Mux.scala 31:69:@2578.4]
  assign _T_5120 = _T_4132 ? 16'h100 : _T_5119; // @[Mux.scala 31:69:@2579.4]
  assign _T_5121 = _T_4129 ? 16'h80 : _T_5120; // @[Mux.scala 31:69:@2580.4]
  assign _T_5122 = _T_4126 ? 16'h40 : _T_5121; // @[Mux.scala 31:69:@2581.4]
  assign _T_5123 = _T_4123 ? 16'h20 : _T_5122; // @[Mux.scala 31:69:@2582.4]
  assign _T_5124 = _T_4168 ? 16'h10 : _T_5123; // @[Mux.scala 31:69:@2583.4]
  assign _T_5125 = _T_4165 ? 16'h8 : _T_5124; // @[Mux.scala 31:69:@2584.4]
  assign _T_5126 = _T_4162 ? 16'h4 : _T_5125; // @[Mux.scala 31:69:@2585.4]
  assign _T_5127 = _T_4159 ? 16'h2 : _T_5126; // @[Mux.scala 31:69:@2586.4]
  assign _T_5128 = _T_4156 ? 16'h1 : _T_5127; // @[Mux.scala 31:69:@2587.4]
  assign _T_5129 = _T_5128[0]; // @[OneHot.scala 66:30:@2588.4]
  assign _T_5130 = _T_5128[1]; // @[OneHot.scala 66:30:@2589.4]
  assign _T_5131 = _T_5128[2]; // @[OneHot.scala 66:30:@2590.4]
  assign _T_5132 = _T_5128[3]; // @[OneHot.scala 66:30:@2591.4]
  assign _T_5133 = _T_5128[4]; // @[OneHot.scala 66:30:@2592.4]
  assign _T_5134 = _T_5128[5]; // @[OneHot.scala 66:30:@2593.4]
  assign _T_5135 = _T_5128[6]; // @[OneHot.scala 66:30:@2594.4]
  assign _T_5136 = _T_5128[7]; // @[OneHot.scala 66:30:@2595.4]
  assign _T_5137 = _T_5128[8]; // @[OneHot.scala 66:30:@2596.4]
  assign _T_5138 = _T_5128[9]; // @[OneHot.scala 66:30:@2597.4]
  assign _T_5139 = _T_5128[10]; // @[OneHot.scala 66:30:@2598.4]
  assign _T_5140 = _T_5128[11]; // @[OneHot.scala 66:30:@2599.4]
  assign _T_5141 = _T_5128[12]; // @[OneHot.scala 66:30:@2600.4]
  assign _T_5142 = _T_5128[13]; // @[OneHot.scala 66:30:@2601.4]
  assign _T_5143 = _T_5128[14]; // @[OneHot.scala 66:30:@2602.4]
  assign _T_5144 = _T_5128[15]; // @[OneHot.scala 66:30:@2603.4]
  assign _T_5185 = _T_4156 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2621.4]
  assign _T_5186 = _T_4153 ? 16'h4000 : _T_5185; // @[Mux.scala 31:69:@2622.4]
  assign _T_5187 = _T_4150 ? 16'h2000 : _T_5186; // @[Mux.scala 31:69:@2623.4]
  assign _T_5188 = _T_4147 ? 16'h1000 : _T_5187; // @[Mux.scala 31:69:@2624.4]
  assign _T_5189 = _T_4144 ? 16'h800 : _T_5188; // @[Mux.scala 31:69:@2625.4]
  assign _T_5190 = _T_4141 ? 16'h400 : _T_5189; // @[Mux.scala 31:69:@2626.4]
  assign _T_5191 = _T_4138 ? 16'h200 : _T_5190; // @[Mux.scala 31:69:@2627.4]
  assign _T_5192 = _T_4135 ? 16'h100 : _T_5191; // @[Mux.scala 31:69:@2628.4]
  assign _T_5193 = _T_4132 ? 16'h80 : _T_5192; // @[Mux.scala 31:69:@2629.4]
  assign _T_5194 = _T_4129 ? 16'h40 : _T_5193; // @[Mux.scala 31:69:@2630.4]
  assign _T_5195 = _T_4126 ? 16'h20 : _T_5194; // @[Mux.scala 31:69:@2631.4]
  assign _T_5196 = _T_4123 ? 16'h10 : _T_5195; // @[Mux.scala 31:69:@2632.4]
  assign _T_5197 = _T_4168 ? 16'h8 : _T_5196; // @[Mux.scala 31:69:@2633.4]
  assign _T_5198 = _T_4165 ? 16'h4 : _T_5197; // @[Mux.scala 31:69:@2634.4]
  assign _T_5199 = _T_4162 ? 16'h2 : _T_5198; // @[Mux.scala 31:69:@2635.4]
  assign _T_5200 = _T_4159 ? 16'h1 : _T_5199; // @[Mux.scala 31:69:@2636.4]
  assign _T_5201 = _T_5200[0]; // @[OneHot.scala 66:30:@2637.4]
  assign _T_5202 = _T_5200[1]; // @[OneHot.scala 66:30:@2638.4]
  assign _T_5203 = _T_5200[2]; // @[OneHot.scala 66:30:@2639.4]
  assign _T_5204 = _T_5200[3]; // @[OneHot.scala 66:30:@2640.4]
  assign _T_5205 = _T_5200[4]; // @[OneHot.scala 66:30:@2641.4]
  assign _T_5206 = _T_5200[5]; // @[OneHot.scala 66:30:@2642.4]
  assign _T_5207 = _T_5200[6]; // @[OneHot.scala 66:30:@2643.4]
  assign _T_5208 = _T_5200[7]; // @[OneHot.scala 66:30:@2644.4]
  assign _T_5209 = _T_5200[8]; // @[OneHot.scala 66:30:@2645.4]
  assign _T_5210 = _T_5200[9]; // @[OneHot.scala 66:30:@2646.4]
  assign _T_5211 = _T_5200[10]; // @[OneHot.scala 66:30:@2647.4]
  assign _T_5212 = _T_5200[11]; // @[OneHot.scala 66:30:@2648.4]
  assign _T_5213 = _T_5200[12]; // @[OneHot.scala 66:30:@2649.4]
  assign _T_5214 = _T_5200[13]; // @[OneHot.scala 66:30:@2650.4]
  assign _T_5215 = _T_5200[14]; // @[OneHot.scala 66:30:@2651.4]
  assign _T_5216 = _T_5200[15]; // @[OneHot.scala 66:30:@2652.4]
  assign _T_5257 = _T_4159 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2670.4]
  assign _T_5258 = _T_4156 ? 16'h4000 : _T_5257; // @[Mux.scala 31:69:@2671.4]
  assign _T_5259 = _T_4153 ? 16'h2000 : _T_5258; // @[Mux.scala 31:69:@2672.4]
  assign _T_5260 = _T_4150 ? 16'h1000 : _T_5259; // @[Mux.scala 31:69:@2673.4]
  assign _T_5261 = _T_4147 ? 16'h800 : _T_5260; // @[Mux.scala 31:69:@2674.4]
  assign _T_5262 = _T_4144 ? 16'h400 : _T_5261; // @[Mux.scala 31:69:@2675.4]
  assign _T_5263 = _T_4141 ? 16'h200 : _T_5262; // @[Mux.scala 31:69:@2676.4]
  assign _T_5264 = _T_4138 ? 16'h100 : _T_5263; // @[Mux.scala 31:69:@2677.4]
  assign _T_5265 = _T_4135 ? 16'h80 : _T_5264; // @[Mux.scala 31:69:@2678.4]
  assign _T_5266 = _T_4132 ? 16'h40 : _T_5265; // @[Mux.scala 31:69:@2679.4]
  assign _T_5267 = _T_4129 ? 16'h20 : _T_5266; // @[Mux.scala 31:69:@2680.4]
  assign _T_5268 = _T_4126 ? 16'h10 : _T_5267; // @[Mux.scala 31:69:@2681.4]
  assign _T_5269 = _T_4123 ? 16'h8 : _T_5268; // @[Mux.scala 31:69:@2682.4]
  assign _T_5270 = _T_4168 ? 16'h4 : _T_5269; // @[Mux.scala 31:69:@2683.4]
  assign _T_5271 = _T_4165 ? 16'h2 : _T_5270; // @[Mux.scala 31:69:@2684.4]
  assign _T_5272 = _T_4162 ? 16'h1 : _T_5271; // @[Mux.scala 31:69:@2685.4]
  assign _T_5273 = _T_5272[0]; // @[OneHot.scala 66:30:@2686.4]
  assign _T_5274 = _T_5272[1]; // @[OneHot.scala 66:30:@2687.4]
  assign _T_5275 = _T_5272[2]; // @[OneHot.scala 66:30:@2688.4]
  assign _T_5276 = _T_5272[3]; // @[OneHot.scala 66:30:@2689.4]
  assign _T_5277 = _T_5272[4]; // @[OneHot.scala 66:30:@2690.4]
  assign _T_5278 = _T_5272[5]; // @[OneHot.scala 66:30:@2691.4]
  assign _T_5279 = _T_5272[6]; // @[OneHot.scala 66:30:@2692.4]
  assign _T_5280 = _T_5272[7]; // @[OneHot.scala 66:30:@2693.4]
  assign _T_5281 = _T_5272[8]; // @[OneHot.scala 66:30:@2694.4]
  assign _T_5282 = _T_5272[9]; // @[OneHot.scala 66:30:@2695.4]
  assign _T_5283 = _T_5272[10]; // @[OneHot.scala 66:30:@2696.4]
  assign _T_5284 = _T_5272[11]; // @[OneHot.scala 66:30:@2697.4]
  assign _T_5285 = _T_5272[12]; // @[OneHot.scala 66:30:@2698.4]
  assign _T_5286 = _T_5272[13]; // @[OneHot.scala 66:30:@2699.4]
  assign _T_5287 = _T_5272[14]; // @[OneHot.scala 66:30:@2700.4]
  assign _T_5288 = _T_5272[15]; // @[OneHot.scala 66:30:@2701.4]
  assign _T_5329 = _T_4162 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2719.4]
  assign _T_5330 = _T_4159 ? 16'h4000 : _T_5329; // @[Mux.scala 31:69:@2720.4]
  assign _T_5331 = _T_4156 ? 16'h2000 : _T_5330; // @[Mux.scala 31:69:@2721.4]
  assign _T_5332 = _T_4153 ? 16'h1000 : _T_5331; // @[Mux.scala 31:69:@2722.4]
  assign _T_5333 = _T_4150 ? 16'h800 : _T_5332; // @[Mux.scala 31:69:@2723.4]
  assign _T_5334 = _T_4147 ? 16'h400 : _T_5333; // @[Mux.scala 31:69:@2724.4]
  assign _T_5335 = _T_4144 ? 16'h200 : _T_5334; // @[Mux.scala 31:69:@2725.4]
  assign _T_5336 = _T_4141 ? 16'h100 : _T_5335; // @[Mux.scala 31:69:@2726.4]
  assign _T_5337 = _T_4138 ? 16'h80 : _T_5336; // @[Mux.scala 31:69:@2727.4]
  assign _T_5338 = _T_4135 ? 16'h40 : _T_5337; // @[Mux.scala 31:69:@2728.4]
  assign _T_5339 = _T_4132 ? 16'h20 : _T_5338; // @[Mux.scala 31:69:@2729.4]
  assign _T_5340 = _T_4129 ? 16'h10 : _T_5339; // @[Mux.scala 31:69:@2730.4]
  assign _T_5341 = _T_4126 ? 16'h8 : _T_5340; // @[Mux.scala 31:69:@2731.4]
  assign _T_5342 = _T_4123 ? 16'h4 : _T_5341; // @[Mux.scala 31:69:@2732.4]
  assign _T_5343 = _T_4168 ? 16'h2 : _T_5342; // @[Mux.scala 31:69:@2733.4]
  assign _T_5344 = _T_4165 ? 16'h1 : _T_5343; // @[Mux.scala 31:69:@2734.4]
  assign _T_5345 = _T_5344[0]; // @[OneHot.scala 66:30:@2735.4]
  assign _T_5346 = _T_5344[1]; // @[OneHot.scala 66:30:@2736.4]
  assign _T_5347 = _T_5344[2]; // @[OneHot.scala 66:30:@2737.4]
  assign _T_5348 = _T_5344[3]; // @[OneHot.scala 66:30:@2738.4]
  assign _T_5349 = _T_5344[4]; // @[OneHot.scala 66:30:@2739.4]
  assign _T_5350 = _T_5344[5]; // @[OneHot.scala 66:30:@2740.4]
  assign _T_5351 = _T_5344[6]; // @[OneHot.scala 66:30:@2741.4]
  assign _T_5352 = _T_5344[7]; // @[OneHot.scala 66:30:@2742.4]
  assign _T_5353 = _T_5344[8]; // @[OneHot.scala 66:30:@2743.4]
  assign _T_5354 = _T_5344[9]; // @[OneHot.scala 66:30:@2744.4]
  assign _T_5355 = _T_5344[10]; // @[OneHot.scala 66:30:@2745.4]
  assign _T_5356 = _T_5344[11]; // @[OneHot.scala 66:30:@2746.4]
  assign _T_5357 = _T_5344[12]; // @[OneHot.scala 66:30:@2747.4]
  assign _T_5358 = _T_5344[13]; // @[OneHot.scala 66:30:@2748.4]
  assign _T_5359 = _T_5344[14]; // @[OneHot.scala 66:30:@2749.4]
  assign _T_5360 = _T_5344[15]; // @[OneHot.scala 66:30:@2750.4]
  assign _T_5401 = _T_4165 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2768.4]
  assign _T_5402 = _T_4162 ? 16'h4000 : _T_5401; // @[Mux.scala 31:69:@2769.4]
  assign _T_5403 = _T_4159 ? 16'h2000 : _T_5402; // @[Mux.scala 31:69:@2770.4]
  assign _T_5404 = _T_4156 ? 16'h1000 : _T_5403; // @[Mux.scala 31:69:@2771.4]
  assign _T_5405 = _T_4153 ? 16'h800 : _T_5404; // @[Mux.scala 31:69:@2772.4]
  assign _T_5406 = _T_4150 ? 16'h400 : _T_5405; // @[Mux.scala 31:69:@2773.4]
  assign _T_5407 = _T_4147 ? 16'h200 : _T_5406; // @[Mux.scala 31:69:@2774.4]
  assign _T_5408 = _T_4144 ? 16'h100 : _T_5407; // @[Mux.scala 31:69:@2775.4]
  assign _T_5409 = _T_4141 ? 16'h80 : _T_5408; // @[Mux.scala 31:69:@2776.4]
  assign _T_5410 = _T_4138 ? 16'h40 : _T_5409; // @[Mux.scala 31:69:@2777.4]
  assign _T_5411 = _T_4135 ? 16'h20 : _T_5410; // @[Mux.scala 31:69:@2778.4]
  assign _T_5412 = _T_4132 ? 16'h10 : _T_5411; // @[Mux.scala 31:69:@2779.4]
  assign _T_5413 = _T_4129 ? 16'h8 : _T_5412; // @[Mux.scala 31:69:@2780.4]
  assign _T_5414 = _T_4126 ? 16'h4 : _T_5413; // @[Mux.scala 31:69:@2781.4]
  assign _T_5415 = _T_4123 ? 16'h2 : _T_5414; // @[Mux.scala 31:69:@2782.4]
  assign _T_5416 = _T_4168 ? 16'h1 : _T_5415; // @[Mux.scala 31:69:@2783.4]
  assign _T_5417 = _T_5416[0]; // @[OneHot.scala 66:30:@2784.4]
  assign _T_5418 = _T_5416[1]; // @[OneHot.scala 66:30:@2785.4]
  assign _T_5419 = _T_5416[2]; // @[OneHot.scala 66:30:@2786.4]
  assign _T_5420 = _T_5416[3]; // @[OneHot.scala 66:30:@2787.4]
  assign _T_5421 = _T_5416[4]; // @[OneHot.scala 66:30:@2788.4]
  assign _T_5422 = _T_5416[5]; // @[OneHot.scala 66:30:@2789.4]
  assign _T_5423 = _T_5416[6]; // @[OneHot.scala 66:30:@2790.4]
  assign _T_5424 = _T_5416[7]; // @[OneHot.scala 66:30:@2791.4]
  assign _T_5425 = _T_5416[8]; // @[OneHot.scala 66:30:@2792.4]
  assign _T_5426 = _T_5416[9]; // @[OneHot.scala 66:30:@2793.4]
  assign _T_5427 = _T_5416[10]; // @[OneHot.scala 66:30:@2794.4]
  assign _T_5428 = _T_5416[11]; // @[OneHot.scala 66:30:@2795.4]
  assign _T_5429 = _T_5416[12]; // @[OneHot.scala 66:30:@2796.4]
  assign _T_5430 = _T_5416[13]; // @[OneHot.scala 66:30:@2797.4]
  assign _T_5431 = _T_5416[14]; // @[OneHot.scala 66:30:@2798.4]
  assign _T_5432 = _T_5416[15]; // @[OneHot.scala 66:30:@2799.4]
  assign _T_5497 = {_T_4344,_T_4343,_T_4342,_T_4341,_T_4340,_T_4339,_T_4338,_T_4337}; // @[Mux.scala 19:72:@2823.4]
  assign _T_5505 = {_T_4352,_T_4351,_T_4350,_T_4349,_T_4348,_T_4347,_T_4346,_T_4345,_T_5497}; // @[Mux.scala 19:72:@2831.4]
  assign _T_5507 = _T_4265 ? _T_5505 : 16'h0; // @[Mux.scala 19:72:@2832.4]
  assign _T_5514 = {_T_4415,_T_4414,_T_4413,_T_4412,_T_4411,_T_4410,_T_4409,_T_4424}; // @[Mux.scala 19:72:@2839.4]
  assign _T_5522 = {_T_4423,_T_4422,_T_4421,_T_4420,_T_4419,_T_4418,_T_4417,_T_4416,_T_5514}; // @[Mux.scala 19:72:@2847.4]
  assign _T_5524 = _T_4266 ? _T_5522 : 16'h0; // @[Mux.scala 19:72:@2848.4]
  assign _T_5531 = {_T_4486,_T_4485,_T_4484,_T_4483,_T_4482,_T_4481,_T_4496,_T_4495}; // @[Mux.scala 19:72:@2855.4]
  assign _T_5539 = {_T_4494,_T_4493,_T_4492,_T_4491,_T_4490,_T_4489,_T_4488,_T_4487,_T_5531}; // @[Mux.scala 19:72:@2863.4]
  assign _T_5541 = _T_4267 ? _T_5539 : 16'h0; // @[Mux.scala 19:72:@2864.4]
  assign _T_5548 = {_T_4557,_T_4556,_T_4555,_T_4554,_T_4553,_T_4568,_T_4567,_T_4566}; // @[Mux.scala 19:72:@2871.4]
  assign _T_5556 = {_T_4565,_T_4564,_T_4563,_T_4562,_T_4561,_T_4560,_T_4559,_T_4558,_T_5548}; // @[Mux.scala 19:72:@2879.4]
  assign _T_5558 = _T_4268 ? _T_5556 : 16'h0; // @[Mux.scala 19:72:@2880.4]
  assign _T_5565 = {_T_4628,_T_4627,_T_4626,_T_4625,_T_4640,_T_4639,_T_4638,_T_4637}; // @[Mux.scala 19:72:@2887.4]
  assign _T_5573 = {_T_4636,_T_4635,_T_4634,_T_4633,_T_4632,_T_4631,_T_4630,_T_4629,_T_5565}; // @[Mux.scala 19:72:@2895.4]
  assign _T_5575 = _T_4269 ? _T_5573 : 16'h0; // @[Mux.scala 19:72:@2896.4]
  assign _T_5582 = {_T_4699,_T_4698,_T_4697,_T_4712,_T_4711,_T_4710,_T_4709,_T_4708}; // @[Mux.scala 19:72:@2903.4]
  assign _T_5590 = {_T_4707,_T_4706,_T_4705,_T_4704,_T_4703,_T_4702,_T_4701,_T_4700,_T_5582}; // @[Mux.scala 19:72:@2911.4]
  assign _T_5592 = _T_4270 ? _T_5590 : 16'h0; // @[Mux.scala 19:72:@2912.4]
  assign _T_5599 = {_T_4770,_T_4769,_T_4784,_T_4783,_T_4782,_T_4781,_T_4780,_T_4779}; // @[Mux.scala 19:72:@2919.4]
  assign _T_5607 = {_T_4778,_T_4777,_T_4776,_T_4775,_T_4774,_T_4773,_T_4772,_T_4771,_T_5599}; // @[Mux.scala 19:72:@2927.4]
  assign _T_5609 = _T_4271 ? _T_5607 : 16'h0; // @[Mux.scala 19:72:@2928.4]
  assign _T_5616 = {_T_4841,_T_4856,_T_4855,_T_4854,_T_4853,_T_4852,_T_4851,_T_4850}; // @[Mux.scala 19:72:@2935.4]
  assign _T_5624 = {_T_4849,_T_4848,_T_4847,_T_4846,_T_4845,_T_4844,_T_4843,_T_4842,_T_5616}; // @[Mux.scala 19:72:@2943.4]
  assign _T_5626 = _T_4272 ? _T_5624 : 16'h0; // @[Mux.scala 19:72:@2944.4]
  assign _T_5633 = {_T_4928,_T_4927,_T_4926,_T_4925,_T_4924,_T_4923,_T_4922,_T_4921}; // @[Mux.scala 19:72:@2951.4]
  assign _T_5641 = {_T_4920,_T_4919,_T_4918,_T_4917,_T_4916,_T_4915,_T_4914,_T_4913,_T_5633}; // @[Mux.scala 19:72:@2959.4]
  assign _T_5643 = _T_4273 ? _T_5641 : 16'h0; // @[Mux.scala 19:72:@2960.4]
  assign _T_5650 = {_T_4999,_T_4998,_T_4997,_T_4996,_T_4995,_T_4994,_T_4993,_T_4992}; // @[Mux.scala 19:72:@2967.4]
  assign _T_5658 = {_T_4991,_T_4990,_T_4989,_T_4988,_T_4987,_T_4986,_T_4985,_T_5000,_T_5650}; // @[Mux.scala 19:72:@2975.4]
  assign _T_5660 = _T_4274 ? _T_5658 : 16'h0; // @[Mux.scala 19:72:@2976.4]
  assign _T_5667 = {_T_5070,_T_5069,_T_5068,_T_5067,_T_5066,_T_5065,_T_5064,_T_5063}; // @[Mux.scala 19:72:@2983.4]
  assign _T_5675 = {_T_5062,_T_5061,_T_5060,_T_5059,_T_5058,_T_5057,_T_5072,_T_5071,_T_5667}; // @[Mux.scala 19:72:@2991.4]
  assign _T_5677 = _T_4275 ? _T_5675 : 16'h0; // @[Mux.scala 19:72:@2992.4]
  assign _T_5684 = {_T_5141,_T_5140,_T_5139,_T_5138,_T_5137,_T_5136,_T_5135,_T_5134}; // @[Mux.scala 19:72:@2999.4]
  assign _T_5692 = {_T_5133,_T_5132,_T_5131,_T_5130,_T_5129,_T_5144,_T_5143,_T_5142,_T_5684}; // @[Mux.scala 19:72:@3007.4]
  assign _T_5694 = _T_4276 ? _T_5692 : 16'h0; // @[Mux.scala 19:72:@3008.4]
  assign _T_5701 = {_T_5212,_T_5211,_T_5210,_T_5209,_T_5208,_T_5207,_T_5206,_T_5205}; // @[Mux.scala 19:72:@3015.4]
  assign _T_5709 = {_T_5204,_T_5203,_T_5202,_T_5201,_T_5216,_T_5215,_T_5214,_T_5213,_T_5701}; // @[Mux.scala 19:72:@3023.4]
  assign _T_5711 = _T_4277 ? _T_5709 : 16'h0; // @[Mux.scala 19:72:@3024.4]
  assign _T_5718 = {_T_5283,_T_5282,_T_5281,_T_5280,_T_5279,_T_5278,_T_5277,_T_5276}; // @[Mux.scala 19:72:@3031.4]
  assign _T_5726 = {_T_5275,_T_5274,_T_5273,_T_5288,_T_5287,_T_5286,_T_5285,_T_5284,_T_5718}; // @[Mux.scala 19:72:@3039.4]
  assign _T_5728 = _T_4278 ? _T_5726 : 16'h0; // @[Mux.scala 19:72:@3040.4]
  assign _T_5735 = {_T_5354,_T_5353,_T_5352,_T_5351,_T_5350,_T_5349,_T_5348,_T_5347}; // @[Mux.scala 19:72:@3047.4]
  assign _T_5743 = {_T_5346,_T_5345,_T_5360,_T_5359,_T_5358,_T_5357,_T_5356,_T_5355,_T_5735}; // @[Mux.scala 19:72:@3055.4]
  assign _T_5745 = _T_4279 ? _T_5743 : 16'h0; // @[Mux.scala 19:72:@3056.4]
  assign _T_5752 = {_T_5425,_T_5424,_T_5423,_T_5422,_T_5421,_T_5420,_T_5419,_T_5418}; // @[Mux.scala 19:72:@3063.4]
  assign _T_5760 = {_T_5417,_T_5432,_T_5431,_T_5430,_T_5429,_T_5428,_T_5427,_T_5426,_T_5752}; // @[Mux.scala 19:72:@3071.4]
  assign _T_5762 = _T_4280 ? _T_5760 : 16'h0; // @[Mux.scala 19:72:@3072.4]
  assign _T_5763 = _T_5507 | _T_5524; // @[Mux.scala 19:72:@3073.4]
  assign _T_5764 = _T_5763 | _T_5541; // @[Mux.scala 19:72:@3074.4]
  assign _T_5765 = _T_5764 | _T_5558; // @[Mux.scala 19:72:@3075.4]
  assign _T_5766 = _T_5765 | _T_5575; // @[Mux.scala 19:72:@3076.4]
  assign _T_5767 = _T_5766 | _T_5592; // @[Mux.scala 19:72:@3077.4]
  assign _T_5768 = _T_5767 | _T_5609; // @[Mux.scala 19:72:@3078.4]
  assign _T_5769 = _T_5768 | _T_5626; // @[Mux.scala 19:72:@3079.4]
  assign _T_5770 = _T_5769 | _T_5643; // @[Mux.scala 19:72:@3080.4]
  assign _T_5771 = _T_5770 | _T_5660; // @[Mux.scala 19:72:@3081.4]
  assign _T_5772 = _T_5771 | _T_5677; // @[Mux.scala 19:72:@3082.4]
  assign _T_5773 = _T_5772 | _T_5694; // @[Mux.scala 19:72:@3083.4]
  assign _T_5774 = _T_5773 | _T_5711; // @[Mux.scala 19:72:@3084.4]
  assign _T_5775 = _T_5774 | _T_5728; // @[Mux.scala 19:72:@3085.4]
  assign _T_5776 = _T_5775 | _T_5745; // @[Mux.scala 19:72:@3086.4]
  assign _T_5777 = _T_5776 | _T_5762; // @[Mux.scala 19:72:@3087.4]
  assign inputAddrPriorityPorts_0_0 = _T_5777[0]; // @[Mux.scala 19:72:@3091.4]
  assign inputAddrPriorityPorts_0_1 = _T_5777[1]; // @[Mux.scala 19:72:@3093.4]
  assign inputAddrPriorityPorts_0_2 = _T_5777[2]; // @[Mux.scala 19:72:@3095.4]
  assign inputAddrPriorityPorts_0_3 = _T_5777[3]; // @[Mux.scala 19:72:@3097.4]
  assign inputAddrPriorityPorts_0_4 = _T_5777[4]; // @[Mux.scala 19:72:@3099.4]
  assign inputAddrPriorityPorts_0_5 = _T_5777[5]; // @[Mux.scala 19:72:@3101.4]
  assign inputAddrPriorityPorts_0_6 = _T_5777[6]; // @[Mux.scala 19:72:@3103.4]
  assign inputAddrPriorityPorts_0_7 = _T_5777[7]; // @[Mux.scala 19:72:@3105.4]
  assign inputAddrPriorityPorts_0_8 = _T_5777[8]; // @[Mux.scala 19:72:@3107.4]
  assign inputAddrPriorityPorts_0_9 = _T_5777[9]; // @[Mux.scala 19:72:@3109.4]
  assign inputAddrPriorityPorts_0_10 = _T_5777[10]; // @[Mux.scala 19:72:@3111.4]
  assign inputAddrPriorityPorts_0_11 = _T_5777[11]; // @[Mux.scala 19:72:@3113.4]
  assign inputAddrPriorityPorts_0_12 = _T_5777[12]; // @[Mux.scala 19:72:@3115.4]
  assign inputAddrPriorityPorts_0_13 = _T_5777[13]; // @[Mux.scala 19:72:@3117.4]
  assign inputAddrPriorityPorts_0_14 = _T_5777[14]; // @[Mux.scala 19:72:@3119.4]
  assign inputAddrPriorityPorts_0_15 = _T_5777[15]; // @[Mux.scala 19:72:@3121.4]
  assign _T_5979 = _T_4238 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3175.4]
  assign _T_5980 = _T_4235 ? 16'h4000 : _T_5979; // @[Mux.scala 31:69:@3176.4]
  assign _T_5981 = _T_4232 ? 16'h2000 : _T_5980; // @[Mux.scala 31:69:@3177.4]
  assign _T_5982 = _T_4229 ? 16'h1000 : _T_5981; // @[Mux.scala 31:69:@3178.4]
  assign _T_5983 = _T_4226 ? 16'h800 : _T_5982; // @[Mux.scala 31:69:@3179.4]
  assign _T_5984 = _T_4223 ? 16'h400 : _T_5983; // @[Mux.scala 31:69:@3180.4]
  assign _T_5985 = _T_4220 ? 16'h200 : _T_5984; // @[Mux.scala 31:69:@3181.4]
  assign _T_5986 = _T_4217 ? 16'h100 : _T_5985; // @[Mux.scala 31:69:@3182.4]
  assign _T_5987 = _T_4214 ? 16'h80 : _T_5986; // @[Mux.scala 31:69:@3183.4]
  assign _T_5988 = _T_4211 ? 16'h40 : _T_5987; // @[Mux.scala 31:69:@3184.4]
  assign _T_5989 = _T_4208 ? 16'h20 : _T_5988; // @[Mux.scala 31:69:@3185.4]
  assign _T_5990 = _T_4205 ? 16'h10 : _T_5989; // @[Mux.scala 31:69:@3186.4]
  assign _T_5991 = _T_4202 ? 16'h8 : _T_5990; // @[Mux.scala 31:69:@3187.4]
  assign _T_5992 = _T_4199 ? 16'h4 : _T_5991; // @[Mux.scala 31:69:@3188.4]
  assign _T_5993 = _T_4196 ? 16'h2 : _T_5992; // @[Mux.scala 31:69:@3189.4]
  assign _T_5994 = _T_4193 ? 16'h1 : _T_5993; // @[Mux.scala 31:69:@3190.4]
  assign _T_5995 = _T_5994[0]; // @[OneHot.scala 66:30:@3191.4]
  assign _T_5996 = _T_5994[1]; // @[OneHot.scala 66:30:@3192.4]
  assign _T_5997 = _T_5994[2]; // @[OneHot.scala 66:30:@3193.4]
  assign _T_5998 = _T_5994[3]; // @[OneHot.scala 66:30:@3194.4]
  assign _T_5999 = _T_5994[4]; // @[OneHot.scala 66:30:@3195.4]
  assign _T_6000 = _T_5994[5]; // @[OneHot.scala 66:30:@3196.4]
  assign _T_6001 = _T_5994[6]; // @[OneHot.scala 66:30:@3197.4]
  assign _T_6002 = _T_5994[7]; // @[OneHot.scala 66:30:@3198.4]
  assign _T_6003 = _T_5994[8]; // @[OneHot.scala 66:30:@3199.4]
  assign _T_6004 = _T_5994[9]; // @[OneHot.scala 66:30:@3200.4]
  assign _T_6005 = _T_5994[10]; // @[OneHot.scala 66:30:@3201.4]
  assign _T_6006 = _T_5994[11]; // @[OneHot.scala 66:30:@3202.4]
  assign _T_6007 = _T_5994[12]; // @[OneHot.scala 66:30:@3203.4]
  assign _T_6008 = _T_5994[13]; // @[OneHot.scala 66:30:@3204.4]
  assign _T_6009 = _T_5994[14]; // @[OneHot.scala 66:30:@3205.4]
  assign _T_6010 = _T_5994[15]; // @[OneHot.scala 66:30:@3206.4]
  assign _T_6051 = _T_4193 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3224.4]
  assign _T_6052 = _T_4238 ? 16'h4000 : _T_6051; // @[Mux.scala 31:69:@3225.4]
  assign _T_6053 = _T_4235 ? 16'h2000 : _T_6052; // @[Mux.scala 31:69:@3226.4]
  assign _T_6054 = _T_4232 ? 16'h1000 : _T_6053; // @[Mux.scala 31:69:@3227.4]
  assign _T_6055 = _T_4229 ? 16'h800 : _T_6054; // @[Mux.scala 31:69:@3228.4]
  assign _T_6056 = _T_4226 ? 16'h400 : _T_6055; // @[Mux.scala 31:69:@3229.4]
  assign _T_6057 = _T_4223 ? 16'h200 : _T_6056; // @[Mux.scala 31:69:@3230.4]
  assign _T_6058 = _T_4220 ? 16'h100 : _T_6057; // @[Mux.scala 31:69:@3231.4]
  assign _T_6059 = _T_4217 ? 16'h80 : _T_6058; // @[Mux.scala 31:69:@3232.4]
  assign _T_6060 = _T_4214 ? 16'h40 : _T_6059; // @[Mux.scala 31:69:@3233.4]
  assign _T_6061 = _T_4211 ? 16'h20 : _T_6060; // @[Mux.scala 31:69:@3234.4]
  assign _T_6062 = _T_4208 ? 16'h10 : _T_6061; // @[Mux.scala 31:69:@3235.4]
  assign _T_6063 = _T_4205 ? 16'h8 : _T_6062; // @[Mux.scala 31:69:@3236.4]
  assign _T_6064 = _T_4202 ? 16'h4 : _T_6063; // @[Mux.scala 31:69:@3237.4]
  assign _T_6065 = _T_4199 ? 16'h2 : _T_6064; // @[Mux.scala 31:69:@3238.4]
  assign _T_6066 = _T_4196 ? 16'h1 : _T_6065; // @[Mux.scala 31:69:@3239.4]
  assign _T_6067 = _T_6066[0]; // @[OneHot.scala 66:30:@3240.4]
  assign _T_6068 = _T_6066[1]; // @[OneHot.scala 66:30:@3241.4]
  assign _T_6069 = _T_6066[2]; // @[OneHot.scala 66:30:@3242.4]
  assign _T_6070 = _T_6066[3]; // @[OneHot.scala 66:30:@3243.4]
  assign _T_6071 = _T_6066[4]; // @[OneHot.scala 66:30:@3244.4]
  assign _T_6072 = _T_6066[5]; // @[OneHot.scala 66:30:@3245.4]
  assign _T_6073 = _T_6066[6]; // @[OneHot.scala 66:30:@3246.4]
  assign _T_6074 = _T_6066[7]; // @[OneHot.scala 66:30:@3247.4]
  assign _T_6075 = _T_6066[8]; // @[OneHot.scala 66:30:@3248.4]
  assign _T_6076 = _T_6066[9]; // @[OneHot.scala 66:30:@3249.4]
  assign _T_6077 = _T_6066[10]; // @[OneHot.scala 66:30:@3250.4]
  assign _T_6078 = _T_6066[11]; // @[OneHot.scala 66:30:@3251.4]
  assign _T_6079 = _T_6066[12]; // @[OneHot.scala 66:30:@3252.4]
  assign _T_6080 = _T_6066[13]; // @[OneHot.scala 66:30:@3253.4]
  assign _T_6081 = _T_6066[14]; // @[OneHot.scala 66:30:@3254.4]
  assign _T_6082 = _T_6066[15]; // @[OneHot.scala 66:30:@3255.4]
  assign _T_6123 = _T_4196 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3273.4]
  assign _T_6124 = _T_4193 ? 16'h4000 : _T_6123; // @[Mux.scala 31:69:@3274.4]
  assign _T_6125 = _T_4238 ? 16'h2000 : _T_6124; // @[Mux.scala 31:69:@3275.4]
  assign _T_6126 = _T_4235 ? 16'h1000 : _T_6125; // @[Mux.scala 31:69:@3276.4]
  assign _T_6127 = _T_4232 ? 16'h800 : _T_6126; // @[Mux.scala 31:69:@3277.4]
  assign _T_6128 = _T_4229 ? 16'h400 : _T_6127; // @[Mux.scala 31:69:@3278.4]
  assign _T_6129 = _T_4226 ? 16'h200 : _T_6128; // @[Mux.scala 31:69:@3279.4]
  assign _T_6130 = _T_4223 ? 16'h100 : _T_6129; // @[Mux.scala 31:69:@3280.4]
  assign _T_6131 = _T_4220 ? 16'h80 : _T_6130; // @[Mux.scala 31:69:@3281.4]
  assign _T_6132 = _T_4217 ? 16'h40 : _T_6131; // @[Mux.scala 31:69:@3282.4]
  assign _T_6133 = _T_4214 ? 16'h20 : _T_6132; // @[Mux.scala 31:69:@3283.4]
  assign _T_6134 = _T_4211 ? 16'h10 : _T_6133; // @[Mux.scala 31:69:@3284.4]
  assign _T_6135 = _T_4208 ? 16'h8 : _T_6134; // @[Mux.scala 31:69:@3285.4]
  assign _T_6136 = _T_4205 ? 16'h4 : _T_6135; // @[Mux.scala 31:69:@3286.4]
  assign _T_6137 = _T_4202 ? 16'h2 : _T_6136; // @[Mux.scala 31:69:@3287.4]
  assign _T_6138 = _T_4199 ? 16'h1 : _T_6137; // @[Mux.scala 31:69:@3288.4]
  assign _T_6139 = _T_6138[0]; // @[OneHot.scala 66:30:@3289.4]
  assign _T_6140 = _T_6138[1]; // @[OneHot.scala 66:30:@3290.4]
  assign _T_6141 = _T_6138[2]; // @[OneHot.scala 66:30:@3291.4]
  assign _T_6142 = _T_6138[3]; // @[OneHot.scala 66:30:@3292.4]
  assign _T_6143 = _T_6138[4]; // @[OneHot.scala 66:30:@3293.4]
  assign _T_6144 = _T_6138[5]; // @[OneHot.scala 66:30:@3294.4]
  assign _T_6145 = _T_6138[6]; // @[OneHot.scala 66:30:@3295.4]
  assign _T_6146 = _T_6138[7]; // @[OneHot.scala 66:30:@3296.4]
  assign _T_6147 = _T_6138[8]; // @[OneHot.scala 66:30:@3297.4]
  assign _T_6148 = _T_6138[9]; // @[OneHot.scala 66:30:@3298.4]
  assign _T_6149 = _T_6138[10]; // @[OneHot.scala 66:30:@3299.4]
  assign _T_6150 = _T_6138[11]; // @[OneHot.scala 66:30:@3300.4]
  assign _T_6151 = _T_6138[12]; // @[OneHot.scala 66:30:@3301.4]
  assign _T_6152 = _T_6138[13]; // @[OneHot.scala 66:30:@3302.4]
  assign _T_6153 = _T_6138[14]; // @[OneHot.scala 66:30:@3303.4]
  assign _T_6154 = _T_6138[15]; // @[OneHot.scala 66:30:@3304.4]
  assign _T_6195 = _T_4199 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3322.4]
  assign _T_6196 = _T_4196 ? 16'h4000 : _T_6195; // @[Mux.scala 31:69:@3323.4]
  assign _T_6197 = _T_4193 ? 16'h2000 : _T_6196; // @[Mux.scala 31:69:@3324.4]
  assign _T_6198 = _T_4238 ? 16'h1000 : _T_6197; // @[Mux.scala 31:69:@3325.4]
  assign _T_6199 = _T_4235 ? 16'h800 : _T_6198; // @[Mux.scala 31:69:@3326.4]
  assign _T_6200 = _T_4232 ? 16'h400 : _T_6199; // @[Mux.scala 31:69:@3327.4]
  assign _T_6201 = _T_4229 ? 16'h200 : _T_6200; // @[Mux.scala 31:69:@3328.4]
  assign _T_6202 = _T_4226 ? 16'h100 : _T_6201; // @[Mux.scala 31:69:@3329.4]
  assign _T_6203 = _T_4223 ? 16'h80 : _T_6202; // @[Mux.scala 31:69:@3330.4]
  assign _T_6204 = _T_4220 ? 16'h40 : _T_6203; // @[Mux.scala 31:69:@3331.4]
  assign _T_6205 = _T_4217 ? 16'h20 : _T_6204; // @[Mux.scala 31:69:@3332.4]
  assign _T_6206 = _T_4214 ? 16'h10 : _T_6205; // @[Mux.scala 31:69:@3333.4]
  assign _T_6207 = _T_4211 ? 16'h8 : _T_6206; // @[Mux.scala 31:69:@3334.4]
  assign _T_6208 = _T_4208 ? 16'h4 : _T_6207; // @[Mux.scala 31:69:@3335.4]
  assign _T_6209 = _T_4205 ? 16'h2 : _T_6208; // @[Mux.scala 31:69:@3336.4]
  assign _T_6210 = _T_4202 ? 16'h1 : _T_6209; // @[Mux.scala 31:69:@3337.4]
  assign _T_6211 = _T_6210[0]; // @[OneHot.scala 66:30:@3338.4]
  assign _T_6212 = _T_6210[1]; // @[OneHot.scala 66:30:@3339.4]
  assign _T_6213 = _T_6210[2]; // @[OneHot.scala 66:30:@3340.4]
  assign _T_6214 = _T_6210[3]; // @[OneHot.scala 66:30:@3341.4]
  assign _T_6215 = _T_6210[4]; // @[OneHot.scala 66:30:@3342.4]
  assign _T_6216 = _T_6210[5]; // @[OneHot.scala 66:30:@3343.4]
  assign _T_6217 = _T_6210[6]; // @[OneHot.scala 66:30:@3344.4]
  assign _T_6218 = _T_6210[7]; // @[OneHot.scala 66:30:@3345.4]
  assign _T_6219 = _T_6210[8]; // @[OneHot.scala 66:30:@3346.4]
  assign _T_6220 = _T_6210[9]; // @[OneHot.scala 66:30:@3347.4]
  assign _T_6221 = _T_6210[10]; // @[OneHot.scala 66:30:@3348.4]
  assign _T_6222 = _T_6210[11]; // @[OneHot.scala 66:30:@3349.4]
  assign _T_6223 = _T_6210[12]; // @[OneHot.scala 66:30:@3350.4]
  assign _T_6224 = _T_6210[13]; // @[OneHot.scala 66:30:@3351.4]
  assign _T_6225 = _T_6210[14]; // @[OneHot.scala 66:30:@3352.4]
  assign _T_6226 = _T_6210[15]; // @[OneHot.scala 66:30:@3353.4]
  assign _T_6267 = _T_4202 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3371.4]
  assign _T_6268 = _T_4199 ? 16'h4000 : _T_6267; // @[Mux.scala 31:69:@3372.4]
  assign _T_6269 = _T_4196 ? 16'h2000 : _T_6268; // @[Mux.scala 31:69:@3373.4]
  assign _T_6270 = _T_4193 ? 16'h1000 : _T_6269; // @[Mux.scala 31:69:@3374.4]
  assign _T_6271 = _T_4238 ? 16'h800 : _T_6270; // @[Mux.scala 31:69:@3375.4]
  assign _T_6272 = _T_4235 ? 16'h400 : _T_6271; // @[Mux.scala 31:69:@3376.4]
  assign _T_6273 = _T_4232 ? 16'h200 : _T_6272; // @[Mux.scala 31:69:@3377.4]
  assign _T_6274 = _T_4229 ? 16'h100 : _T_6273; // @[Mux.scala 31:69:@3378.4]
  assign _T_6275 = _T_4226 ? 16'h80 : _T_6274; // @[Mux.scala 31:69:@3379.4]
  assign _T_6276 = _T_4223 ? 16'h40 : _T_6275; // @[Mux.scala 31:69:@3380.4]
  assign _T_6277 = _T_4220 ? 16'h20 : _T_6276; // @[Mux.scala 31:69:@3381.4]
  assign _T_6278 = _T_4217 ? 16'h10 : _T_6277; // @[Mux.scala 31:69:@3382.4]
  assign _T_6279 = _T_4214 ? 16'h8 : _T_6278; // @[Mux.scala 31:69:@3383.4]
  assign _T_6280 = _T_4211 ? 16'h4 : _T_6279; // @[Mux.scala 31:69:@3384.4]
  assign _T_6281 = _T_4208 ? 16'h2 : _T_6280; // @[Mux.scala 31:69:@3385.4]
  assign _T_6282 = _T_4205 ? 16'h1 : _T_6281; // @[Mux.scala 31:69:@3386.4]
  assign _T_6283 = _T_6282[0]; // @[OneHot.scala 66:30:@3387.4]
  assign _T_6284 = _T_6282[1]; // @[OneHot.scala 66:30:@3388.4]
  assign _T_6285 = _T_6282[2]; // @[OneHot.scala 66:30:@3389.4]
  assign _T_6286 = _T_6282[3]; // @[OneHot.scala 66:30:@3390.4]
  assign _T_6287 = _T_6282[4]; // @[OneHot.scala 66:30:@3391.4]
  assign _T_6288 = _T_6282[5]; // @[OneHot.scala 66:30:@3392.4]
  assign _T_6289 = _T_6282[6]; // @[OneHot.scala 66:30:@3393.4]
  assign _T_6290 = _T_6282[7]; // @[OneHot.scala 66:30:@3394.4]
  assign _T_6291 = _T_6282[8]; // @[OneHot.scala 66:30:@3395.4]
  assign _T_6292 = _T_6282[9]; // @[OneHot.scala 66:30:@3396.4]
  assign _T_6293 = _T_6282[10]; // @[OneHot.scala 66:30:@3397.4]
  assign _T_6294 = _T_6282[11]; // @[OneHot.scala 66:30:@3398.4]
  assign _T_6295 = _T_6282[12]; // @[OneHot.scala 66:30:@3399.4]
  assign _T_6296 = _T_6282[13]; // @[OneHot.scala 66:30:@3400.4]
  assign _T_6297 = _T_6282[14]; // @[OneHot.scala 66:30:@3401.4]
  assign _T_6298 = _T_6282[15]; // @[OneHot.scala 66:30:@3402.4]
  assign _T_6339 = _T_4205 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3420.4]
  assign _T_6340 = _T_4202 ? 16'h4000 : _T_6339; // @[Mux.scala 31:69:@3421.4]
  assign _T_6341 = _T_4199 ? 16'h2000 : _T_6340; // @[Mux.scala 31:69:@3422.4]
  assign _T_6342 = _T_4196 ? 16'h1000 : _T_6341; // @[Mux.scala 31:69:@3423.4]
  assign _T_6343 = _T_4193 ? 16'h800 : _T_6342; // @[Mux.scala 31:69:@3424.4]
  assign _T_6344 = _T_4238 ? 16'h400 : _T_6343; // @[Mux.scala 31:69:@3425.4]
  assign _T_6345 = _T_4235 ? 16'h200 : _T_6344; // @[Mux.scala 31:69:@3426.4]
  assign _T_6346 = _T_4232 ? 16'h100 : _T_6345; // @[Mux.scala 31:69:@3427.4]
  assign _T_6347 = _T_4229 ? 16'h80 : _T_6346; // @[Mux.scala 31:69:@3428.4]
  assign _T_6348 = _T_4226 ? 16'h40 : _T_6347; // @[Mux.scala 31:69:@3429.4]
  assign _T_6349 = _T_4223 ? 16'h20 : _T_6348; // @[Mux.scala 31:69:@3430.4]
  assign _T_6350 = _T_4220 ? 16'h10 : _T_6349; // @[Mux.scala 31:69:@3431.4]
  assign _T_6351 = _T_4217 ? 16'h8 : _T_6350; // @[Mux.scala 31:69:@3432.4]
  assign _T_6352 = _T_4214 ? 16'h4 : _T_6351; // @[Mux.scala 31:69:@3433.4]
  assign _T_6353 = _T_4211 ? 16'h2 : _T_6352; // @[Mux.scala 31:69:@3434.4]
  assign _T_6354 = _T_4208 ? 16'h1 : _T_6353; // @[Mux.scala 31:69:@3435.4]
  assign _T_6355 = _T_6354[0]; // @[OneHot.scala 66:30:@3436.4]
  assign _T_6356 = _T_6354[1]; // @[OneHot.scala 66:30:@3437.4]
  assign _T_6357 = _T_6354[2]; // @[OneHot.scala 66:30:@3438.4]
  assign _T_6358 = _T_6354[3]; // @[OneHot.scala 66:30:@3439.4]
  assign _T_6359 = _T_6354[4]; // @[OneHot.scala 66:30:@3440.4]
  assign _T_6360 = _T_6354[5]; // @[OneHot.scala 66:30:@3441.4]
  assign _T_6361 = _T_6354[6]; // @[OneHot.scala 66:30:@3442.4]
  assign _T_6362 = _T_6354[7]; // @[OneHot.scala 66:30:@3443.4]
  assign _T_6363 = _T_6354[8]; // @[OneHot.scala 66:30:@3444.4]
  assign _T_6364 = _T_6354[9]; // @[OneHot.scala 66:30:@3445.4]
  assign _T_6365 = _T_6354[10]; // @[OneHot.scala 66:30:@3446.4]
  assign _T_6366 = _T_6354[11]; // @[OneHot.scala 66:30:@3447.4]
  assign _T_6367 = _T_6354[12]; // @[OneHot.scala 66:30:@3448.4]
  assign _T_6368 = _T_6354[13]; // @[OneHot.scala 66:30:@3449.4]
  assign _T_6369 = _T_6354[14]; // @[OneHot.scala 66:30:@3450.4]
  assign _T_6370 = _T_6354[15]; // @[OneHot.scala 66:30:@3451.4]
  assign _T_6411 = _T_4208 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3469.4]
  assign _T_6412 = _T_4205 ? 16'h4000 : _T_6411; // @[Mux.scala 31:69:@3470.4]
  assign _T_6413 = _T_4202 ? 16'h2000 : _T_6412; // @[Mux.scala 31:69:@3471.4]
  assign _T_6414 = _T_4199 ? 16'h1000 : _T_6413; // @[Mux.scala 31:69:@3472.4]
  assign _T_6415 = _T_4196 ? 16'h800 : _T_6414; // @[Mux.scala 31:69:@3473.4]
  assign _T_6416 = _T_4193 ? 16'h400 : _T_6415; // @[Mux.scala 31:69:@3474.4]
  assign _T_6417 = _T_4238 ? 16'h200 : _T_6416; // @[Mux.scala 31:69:@3475.4]
  assign _T_6418 = _T_4235 ? 16'h100 : _T_6417; // @[Mux.scala 31:69:@3476.4]
  assign _T_6419 = _T_4232 ? 16'h80 : _T_6418; // @[Mux.scala 31:69:@3477.4]
  assign _T_6420 = _T_4229 ? 16'h40 : _T_6419; // @[Mux.scala 31:69:@3478.4]
  assign _T_6421 = _T_4226 ? 16'h20 : _T_6420; // @[Mux.scala 31:69:@3479.4]
  assign _T_6422 = _T_4223 ? 16'h10 : _T_6421; // @[Mux.scala 31:69:@3480.4]
  assign _T_6423 = _T_4220 ? 16'h8 : _T_6422; // @[Mux.scala 31:69:@3481.4]
  assign _T_6424 = _T_4217 ? 16'h4 : _T_6423; // @[Mux.scala 31:69:@3482.4]
  assign _T_6425 = _T_4214 ? 16'h2 : _T_6424; // @[Mux.scala 31:69:@3483.4]
  assign _T_6426 = _T_4211 ? 16'h1 : _T_6425; // @[Mux.scala 31:69:@3484.4]
  assign _T_6427 = _T_6426[0]; // @[OneHot.scala 66:30:@3485.4]
  assign _T_6428 = _T_6426[1]; // @[OneHot.scala 66:30:@3486.4]
  assign _T_6429 = _T_6426[2]; // @[OneHot.scala 66:30:@3487.4]
  assign _T_6430 = _T_6426[3]; // @[OneHot.scala 66:30:@3488.4]
  assign _T_6431 = _T_6426[4]; // @[OneHot.scala 66:30:@3489.4]
  assign _T_6432 = _T_6426[5]; // @[OneHot.scala 66:30:@3490.4]
  assign _T_6433 = _T_6426[6]; // @[OneHot.scala 66:30:@3491.4]
  assign _T_6434 = _T_6426[7]; // @[OneHot.scala 66:30:@3492.4]
  assign _T_6435 = _T_6426[8]; // @[OneHot.scala 66:30:@3493.4]
  assign _T_6436 = _T_6426[9]; // @[OneHot.scala 66:30:@3494.4]
  assign _T_6437 = _T_6426[10]; // @[OneHot.scala 66:30:@3495.4]
  assign _T_6438 = _T_6426[11]; // @[OneHot.scala 66:30:@3496.4]
  assign _T_6439 = _T_6426[12]; // @[OneHot.scala 66:30:@3497.4]
  assign _T_6440 = _T_6426[13]; // @[OneHot.scala 66:30:@3498.4]
  assign _T_6441 = _T_6426[14]; // @[OneHot.scala 66:30:@3499.4]
  assign _T_6442 = _T_6426[15]; // @[OneHot.scala 66:30:@3500.4]
  assign _T_6483 = _T_4211 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3518.4]
  assign _T_6484 = _T_4208 ? 16'h4000 : _T_6483; // @[Mux.scala 31:69:@3519.4]
  assign _T_6485 = _T_4205 ? 16'h2000 : _T_6484; // @[Mux.scala 31:69:@3520.4]
  assign _T_6486 = _T_4202 ? 16'h1000 : _T_6485; // @[Mux.scala 31:69:@3521.4]
  assign _T_6487 = _T_4199 ? 16'h800 : _T_6486; // @[Mux.scala 31:69:@3522.4]
  assign _T_6488 = _T_4196 ? 16'h400 : _T_6487; // @[Mux.scala 31:69:@3523.4]
  assign _T_6489 = _T_4193 ? 16'h200 : _T_6488; // @[Mux.scala 31:69:@3524.4]
  assign _T_6490 = _T_4238 ? 16'h100 : _T_6489; // @[Mux.scala 31:69:@3525.4]
  assign _T_6491 = _T_4235 ? 16'h80 : _T_6490; // @[Mux.scala 31:69:@3526.4]
  assign _T_6492 = _T_4232 ? 16'h40 : _T_6491; // @[Mux.scala 31:69:@3527.4]
  assign _T_6493 = _T_4229 ? 16'h20 : _T_6492; // @[Mux.scala 31:69:@3528.4]
  assign _T_6494 = _T_4226 ? 16'h10 : _T_6493; // @[Mux.scala 31:69:@3529.4]
  assign _T_6495 = _T_4223 ? 16'h8 : _T_6494; // @[Mux.scala 31:69:@3530.4]
  assign _T_6496 = _T_4220 ? 16'h4 : _T_6495; // @[Mux.scala 31:69:@3531.4]
  assign _T_6497 = _T_4217 ? 16'h2 : _T_6496; // @[Mux.scala 31:69:@3532.4]
  assign _T_6498 = _T_4214 ? 16'h1 : _T_6497; // @[Mux.scala 31:69:@3533.4]
  assign _T_6499 = _T_6498[0]; // @[OneHot.scala 66:30:@3534.4]
  assign _T_6500 = _T_6498[1]; // @[OneHot.scala 66:30:@3535.4]
  assign _T_6501 = _T_6498[2]; // @[OneHot.scala 66:30:@3536.4]
  assign _T_6502 = _T_6498[3]; // @[OneHot.scala 66:30:@3537.4]
  assign _T_6503 = _T_6498[4]; // @[OneHot.scala 66:30:@3538.4]
  assign _T_6504 = _T_6498[5]; // @[OneHot.scala 66:30:@3539.4]
  assign _T_6505 = _T_6498[6]; // @[OneHot.scala 66:30:@3540.4]
  assign _T_6506 = _T_6498[7]; // @[OneHot.scala 66:30:@3541.4]
  assign _T_6507 = _T_6498[8]; // @[OneHot.scala 66:30:@3542.4]
  assign _T_6508 = _T_6498[9]; // @[OneHot.scala 66:30:@3543.4]
  assign _T_6509 = _T_6498[10]; // @[OneHot.scala 66:30:@3544.4]
  assign _T_6510 = _T_6498[11]; // @[OneHot.scala 66:30:@3545.4]
  assign _T_6511 = _T_6498[12]; // @[OneHot.scala 66:30:@3546.4]
  assign _T_6512 = _T_6498[13]; // @[OneHot.scala 66:30:@3547.4]
  assign _T_6513 = _T_6498[14]; // @[OneHot.scala 66:30:@3548.4]
  assign _T_6514 = _T_6498[15]; // @[OneHot.scala 66:30:@3549.4]
  assign _T_6555 = _T_4214 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3567.4]
  assign _T_6556 = _T_4211 ? 16'h4000 : _T_6555; // @[Mux.scala 31:69:@3568.4]
  assign _T_6557 = _T_4208 ? 16'h2000 : _T_6556; // @[Mux.scala 31:69:@3569.4]
  assign _T_6558 = _T_4205 ? 16'h1000 : _T_6557; // @[Mux.scala 31:69:@3570.4]
  assign _T_6559 = _T_4202 ? 16'h800 : _T_6558; // @[Mux.scala 31:69:@3571.4]
  assign _T_6560 = _T_4199 ? 16'h400 : _T_6559; // @[Mux.scala 31:69:@3572.4]
  assign _T_6561 = _T_4196 ? 16'h200 : _T_6560; // @[Mux.scala 31:69:@3573.4]
  assign _T_6562 = _T_4193 ? 16'h100 : _T_6561; // @[Mux.scala 31:69:@3574.4]
  assign _T_6563 = _T_4238 ? 16'h80 : _T_6562; // @[Mux.scala 31:69:@3575.4]
  assign _T_6564 = _T_4235 ? 16'h40 : _T_6563; // @[Mux.scala 31:69:@3576.4]
  assign _T_6565 = _T_4232 ? 16'h20 : _T_6564; // @[Mux.scala 31:69:@3577.4]
  assign _T_6566 = _T_4229 ? 16'h10 : _T_6565; // @[Mux.scala 31:69:@3578.4]
  assign _T_6567 = _T_4226 ? 16'h8 : _T_6566; // @[Mux.scala 31:69:@3579.4]
  assign _T_6568 = _T_4223 ? 16'h4 : _T_6567; // @[Mux.scala 31:69:@3580.4]
  assign _T_6569 = _T_4220 ? 16'h2 : _T_6568; // @[Mux.scala 31:69:@3581.4]
  assign _T_6570 = _T_4217 ? 16'h1 : _T_6569; // @[Mux.scala 31:69:@3582.4]
  assign _T_6571 = _T_6570[0]; // @[OneHot.scala 66:30:@3583.4]
  assign _T_6572 = _T_6570[1]; // @[OneHot.scala 66:30:@3584.4]
  assign _T_6573 = _T_6570[2]; // @[OneHot.scala 66:30:@3585.4]
  assign _T_6574 = _T_6570[3]; // @[OneHot.scala 66:30:@3586.4]
  assign _T_6575 = _T_6570[4]; // @[OneHot.scala 66:30:@3587.4]
  assign _T_6576 = _T_6570[5]; // @[OneHot.scala 66:30:@3588.4]
  assign _T_6577 = _T_6570[6]; // @[OneHot.scala 66:30:@3589.4]
  assign _T_6578 = _T_6570[7]; // @[OneHot.scala 66:30:@3590.4]
  assign _T_6579 = _T_6570[8]; // @[OneHot.scala 66:30:@3591.4]
  assign _T_6580 = _T_6570[9]; // @[OneHot.scala 66:30:@3592.4]
  assign _T_6581 = _T_6570[10]; // @[OneHot.scala 66:30:@3593.4]
  assign _T_6582 = _T_6570[11]; // @[OneHot.scala 66:30:@3594.4]
  assign _T_6583 = _T_6570[12]; // @[OneHot.scala 66:30:@3595.4]
  assign _T_6584 = _T_6570[13]; // @[OneHot.scala 66:30:@3596.4]
  assign _T_6585 = _T_6570[14]; // @[OneHot.scala 66:30:@3597.4]
  assign _T_6586 = _T_6570[15]; // @[OneHot.scala 66:30:@3598.4]
  assign _T_6627 = _T_4217 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3616.4]
  assign _T_6628 = _T_4214 ? 16'h4000 : _T_6627; // @[Mux.scala 31:69:@3617.4]
  assign _T_6629 = _T_4211 ? 16'h2000 : _T_6628; // @[Mux.scala 31:69:@3618.4]
  assign _T_6630 = _T_4208 ? 16'h1000 : _T_6629; // @[Mux.scala 31:69:@3619.4]
  assign _T_6631 = _T_4205 ? 16'h800 : _T_6630; // @[Mux.scala 31:69:@3620.4]
  assign _T_6632 = _T_4202 ? 16'h400 : _T_6631; // @[Mux.scala 31:69:@3621.4]
  assign _T_6633 = _T_4199 ? 16'h200 : _T_6632; // @[Mux.scala 31:69:@3622.4]
  assign _T_6634 = _T_4196 ? 16'h100 : _T_6633; // @[Mux.scala 31:69:@3623.4]
  assign _T_6635 = _T_4193 ? 16'h80 : _T_6634; // @[Mux.scala 31:69:@3624.4]
  assign _T_6636 = _T_4238 ? 16'h40 : _T_6635; // @[Mux.scala 31:69:@3625.4]
  assign _T_6637 = _T_4235 ? 16'h20 : _T_6636; // @[Mux.scala 31:69:@3626.4]
  assign _T_6638 = _T_4232 ? 16'h10 : _T_6637; // @[Mux.scala 31:69:@3627.4]
  assign _T_6639 = _T_4229 ? 16'h8 : _T_6638; // @[Mux.scala 31:69:@3628.4]
  assign _T_6640 = _T_4226 ? 16'h4 : _T_6639; // @[Mux.scala 31:69:@3629.4]
  assign _T_6641 = _T_4223 ? 16'h2 : _T_6640; // @[Mux.scala 31:69:@3630.4]
  assign _T_6642 = _T_4220 ? 16'h1 : _T_6641; // @[Mux.scala 31:69:@3631.4]
  assign _T_6643 = _T_6642[0]; // @[OneHot.scala 66:30:@3632.4]
  assign _T_6644 = _T_6642[1]; // @[OneHot.scala 66:30:@3633.4]
  assign _T_6645 = _T_6642[2]; // @[OneHot.scala 66:30:@3634.4]
  assign _T_6646 = _T_6642[3]; // @[OneHot.scala 66:30:@3635.4]
  assign _T_6647 = _T_6642[4]; // @[OneHot.scala 66:30:@3636.4]
  assign _T_6648 = _T_6642[5]; // @[OneHot.scala 66:30:@3637.4]
  assign _T_6649 = _T_6642[6]; // @[OneHot.scala 66:30:@3638.4]
  assign _T_6650 = _T_6642[7]; // @[OneHot.scala 66:30:@3639.4]
  assign _T_6651 = _T_6642[8]; // @[OneHot.scala 66:30:@3640.4]
  assign _T_6652 = _T_6642[9]; // @[OneHot.scala 66:30:@3641.4]
  assign _T_6653 = _T_6642[10]; // @[OneHot.scala 66:30:@3642.4]
  assign _T_6654 = _T_6642[11]; // @[OneHot.scala 66:30:@3643.4]
  assign _T_6655 = _T_6642[12]; // @[OneHot.scala 66:30:@3644.4]
  assign _T_6656 = _T_6642[13]; // @[OneHot.scala 66:30:@3645.4]
  assign _T_6657 = _T_6642[14]; // @[OneHot.scala 66:30:@3646.4]
  assign _T_6658 = _T_6642[15]; // @[OneHot.scala 66:30:@3647.4]
  assign _T_6699 = _T_4220 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3665.4]
  assign _T_6700 = _T_4217 ? 16'h4000 : _T_6699; // @[Mux.scala 31:69:@3666.4]
  assign _T_6701 = _T_4214 ? 16'h2000 : _T_6700; // @[Mux.scala 31:69:@3667.4]
  assign _T_6702 = _T_4211 ? 16'h1000 : _T_6701; // @[Mux.scala 31:69:@3668.4]
  assign _T_6703 = _T_4208 ? 16'h800 : _T_6702; // @[Mux.scala 31:69:@3669.4]
  assign _T_6704 = _T_4205 ? 16'h400 : _T_6703; // @[Mux.scala 31:69:@3670.4]
  assign _T_6705 = _T_4202 ? 16'h200 : _T_6704; // @[Mux.scala 31:69:@3671.4]
  assign _T_6706 = _T_4199 ? 16'h100 : _T_6705; // @[Mux.scala 31:69:@3672.4]
  assign _T_6707 = _T_4196 ? 16'h80 : _T_6706; // @[Mux.scala 31:69:@3673.4]
  assign _T_6708 = _T_4193 ? 16'h40 : _T_6707; // @[Mux.scala 31:69:@3674.4]
  assign _T_6709 = _T_4238 ? 16'h20 : _T_6708; // @[Mux.scala 31:69:@3675.4]
  assign _T_6710 = _T_4235 ? 16'h10 : _T_6709; // @[Mux.scala 31:69:@3676.4]
  assign _T_6711 = _T_4232 ? 16'h8 : _T_6710; // @[Mux.scala 31:69:@3677.4]
  assign _T_6712 = _T_4229 ? 16'h4 : _T_6711; // @[Mux.scala 31:69:@3678.4]
  assign _T_6713 = _T_4226 ? 16'h2 : _T_6712; // @[Mux.scala 31:69:@3679.4]
  assign _T_6714 = _T_4223 ? 16'h1 : _T_6713; // @[Mux.scala 31:69:@3680.4]
  assign _T_6715 = _T_6714[0]; // @[OneHot.scala 66:30:@3681.4]
  assign _T_6716 = _T_6714[1]; // @[OneHot.scala 66:30:@3682.4]
  assign _T_6717 = _T_6714[2]; // @[OneHot.scala 66:30:@3683.4]
  assign _T_6718 = _T_6714[3]; // @[OneHot.scala 66:30:@3684.4]
  assign _T_6719 = _T_6714[4]; // @[OneHot.scala 66:30:@3685.4]
  assign _T_6720 = _T_6714[5]; // @[OneHot.scala 66:30:@3686.4]
  assign _T_6721 = _T_6714[6]; // @[OneHot.scala 66:30:@3687.4]
  assign _T_6722 = _T_6714[7]; // @[OneHot.scala 66:30:@3688.4]
  assign _T_6723 = _T_6714[8]; // @[OneHot.scala 66:30:@3689.4]
  assign _T_6724 = _T_6714[9]; // @[OneHot.scala 66:30:@3690.4]
  assign _T_6725 = _T_6714[10]; // @[OneHot.scala 66:30:@3691.4]
  assign _T_6726 = _T_6714[11]; // @[OneHot.scala 66:30:@3692.4]
  assign _T_6727 = _T_6714[12]; // @[OneHot.scala 66:30:@3693.4]
  assign _T_6728 = _T_6714[13]; // @[OneHot.scala 66:30:@3694.4]
  assign _T_6729 = _T_6714[14]; // @[OneHot.scala 66:30:@3695.4]
  assign _T_6730 = _T_6714[15]; // @[OneHot.scala 66:30:@3696.4]
  assign _T_6771 = _T_4223 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3714.4]
  assign _T_6772 = _T_4220 ? 16'h4000 : _T_6771; // @[Mux.scala 31:69:@3715.4]
  assign _T_6773 = _T_4217 ? 16'h2000 : _T_6772; // @[Mux.scala 31:69:@3716.4]
  assign _T_6774 = _T_4214 ? 16'h1000 : _T_6773; // @[Mux.scala 31:69:@3717.4]
  assign _T_6775 = _T_4211 ? 16'h800 : _T_6774; // @[Mux.scala 31:69:@3718.4]
  assign _T_6776 = _T_4208 ? 16'h400 : _T_6775; // @[Mux.scala 31:69:@3719.4]
  assign _T_6777 = _T_4205 ? 16'h200 : _T_6776; // @[Mux.scala 31:69:@3720.4]
  assign _T_6778 = _T_4202 ? 16'h100 : _T_6777; // @[Mux.scala 31:69:@3721.4]
  assign _T_6779 = _T_4199 ? 16'h80 : _T_6778; // @[Mux.scala 31:69:@3722.4]
  assign _T_6780 = _T_4196 ? 16'h40 : _T_6779; // @[Mux.scala 31:69:@3723.4]
  assign _T_6781 = _T_4193 ? 16'h20 : _T_6780; // @[Mux.scala 31:69:@3724.4]
  assign _T_6782 = _T_4238 ? 16'h10 : _T_6781; // @[Mux.scala 31:69:@3725.4]
  assign _T_6783 = _T_4235 ? 16'h8 : _T_6782; // @[Mux.scala 31:69:@3726.4]
  assign _T_6784 = _T_4232 ? 16'h4 : _T_6783; // @[Mux.scala 31:69:@3727.4]
  assign _T_6785 = _T_4229 ? 16'h2 : _T_6784; // @[Mux.scala 31:69:@3728.4]
  assign _T_6786 = _T_4226 ? 16'h1 : _T_6785; // @[Mux.scala 31:69:@3729.4]
  assign _T_6787 = _T_6786[0]; // @[OneHot.scala 66:30:@3730.4]
  assign _T_6788 = _T_6786[1]; // @[OneHot.scala 66:30:@3731.4]
  assign _T_6789 = _T_6786[2]; // @[OneHot.scala 66:30:@3732.4]
  assign _T_6790 = _T_6786[3]; // @[OneHot.scala 66:30:@3733.4]
  assign _T_6791 = _T_6786[4]; // @[OneHot.scala 66:30:@3734.4]
  assign _T_6792 = _T_6786[5]; // @[OneHot.scala 66:30:@3735.4]
  assign _T_6793 = _T_6786[6]; // @[OneHot.scala 66:30:@3736.4]
  assign _T_6794 = _T_6786[7]; // @[OneHot.scala 66:30:@3737.4]
  assign _T_6795 = _T_6786[8]; // @[OneHot.scala 66:30:@3738.4]
  assign _T_6796 = _T_6786[9]; // @[OneHot.scala 66:30:@3739.4]
  assign _T_6797 = _T_6786[10]; // @[OneHot.scala 66:30:@3740.4]
  assign _T_6798 = _T_6786[11]; // @[OneHot.scala 66:30:@3741.4]
  assign _T_6799 = _T_6786[12]; // @[OneHot.scala 66:30:@3742.4]
  assign _T_6800 = _T_6786[13]; // @[OneHot.scala 66:30:@3743.4]
  assign _T_6801 = _T_6786[14]; // @[OneHot.scala 66:30:@3744.4]
  assign _T_6802 = _T_6786[15]; // @[OneHot.scala 66:30:@3745.4]
  assign _T_6843 = _T_4226 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3763.4]
  assign _T_6844 = _T_4223 ? 16'h4000 : _T_6843; // @[Mux.scala 31:69:@3764.4]
  assign _T_6845 = _T_4220 ? 16'h2000 : _T_6844; // @[Mux.scala 31:69:@3765.4]
  assign _T_6846 = _T_4217 ? 16'h1000 : _T_6845; // @[Mux.scala 31:69:@3766.4]
  assign _T_6847 = _T_4214 ? 16'h800 : _T_6846; // @[Mux.scala 31:69:@3767.4]
  assign _T_6848 = _T_4211 ? 16'h400 : _T_6847; // @[Mux.scala 31:69:@3768.4]
  assign _T_6849 = _T_4208 ? 16'h200 : _T_6848; // @[Mux.scala 31:69:@3769.4]
  assign _T_6850 = _T_4205 ? 16'h100 : _T_6849; // @[Mux.scala 31:69:@3770.4]
  assign _T_6851 = _T_4202 ? 16'h80 : _T_6850; // @[Mux.scala 31:69:@3771.4]
  assign _T_6852 = _T_4199 ? 16'h40 : _T_6851; // @[Mux.scala 31:69:@3772.4]
  assign _T_6853 = _T_4196 ? 16'h20 : _T_6852; // @[Mux.scala 31:69:@3773.4]
  assign _T_6854 = _T_4193 ? 16'h10 : _T_6853; // @[Mux.scala 31:69:@3774.4]
  assign _T_6855 = _T_4238 ? 16'h8 : _T_6854; // @[Mux.scala 31:69:@3775.4]
  assign _T_6856 = _T_4235 ? 16'h4 : _T_6855; // @[Mux.scala 31:69:@3776.4]
  assign _T_6857 = _T_4232 ? 16'h2 : _T_6856; // @[Mux.scala 31:69:@3777.4]
  assign _T_6858 = _T_4229 ? 16'h1 : _T_6857; // @[Mux.scala 31:69:@3778.4]
  assign _T_6859 = _T_6858[0]; // @[OneHot.scala 66:30:@3779.4]
  assign _T_6860 = _T_6858[1]; // @[OneHot.scala 66:30:@3780.4]
  assign _T_6861 = _T_6858[2]; // @[OneHot.scala 66:30:@3781.4]
  assign _T_6862 = _T_6858[3]; // @[OneHot.scala 66:30:@3782.4]
  assign _T_6863 = _T_6858[4]; // @[OneHot.scala 66:30:@3783.4]
  assign _T_6864 = _T_6858[5]; // @[OneHot.scala 66:30:@3784.4]
  assign _T_6865 = _T_6858[6]; // @[OneHot.scala 66:30:@3785.4]
  assign _T_6866 = _T_6858[7]; // @[OneHot.scala 66:30:@3786.4]
  assign _T_6867 = _T_6858[8]; // @[OneHot.scala 66:30:@3787.4]
  assign _T_6868 = _T_6858[9]; // @[OneHot.scala 66:30:@3788.4]
  assign _T_6869 = _T_6858[10]; // @[OneHot.scala 66:30:@3789.4]
  assign _T_6870 = _T_6858[11]; // @[OneHot.scala 66:30:@3790.4]
  assign _T_6871 = _T_6858[12]; // @[OneHot.scala 66:30:@3791.4]
  assign _T_6872 = _T_6858[13]; // @[OneHot.scala 66:30:@3792.4]
  assign _T_6873 = _T_6858[14]; // @[OneHot.scala 66:30:@3793.4]
  assign _T_6874 = _T_6858[15]; // @[OneHot.scala 66:30:@3794.4]
  assign _T_6915 = _T_4229 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3812.4]
  assign _T_6916 = _T_4226 ? 16'h4000 : _T_6915; // @[Mux.scala 31:69:@3813.4]
  assign _T_6917 = _T_4223 ? 16'h2000 : _T_6916; // @[Mux.scala 31:69:@3814.4]
  assign _T_6918 = _T_4220 ? 16'h1000 : _T_6917; // @[Mux.scala 31:69:@3815.4]
  assign _T_6919 = _T_4217 ? 16'h800 : _T_6918; // @[Mux.scala 31:69:@3816.4]
  assign _T_6920 = _T_4214 ? 16'h400 : _T_6919; // @[Mux.scala 31:69:@3817.4]
  assign _T_6921 = _T_4211 ? 16'h200 : _T_6920; // @[Mux.scala 31:69:@3818.4]
  assign _T_6922 = _T_4208 ? 16'h100 : _T_6921; // @[Mux.scala 31:69:@3819.4]
  assign _T_6923 = _T_4205 ? 16'h80 : _T_6922; // @[Mux.scala 31:69:@3820.4]
  assign _T_6924 = _T_4202 ? 16'h40 : _T_6923; // @[Mux.scala 31:69:@3821.4]
  assign _T_6925 = _T_4199 ? 16'h20 : _T_6924; // @[Mux.scala 31:69:@3822.4]
  assign _T_6926 = _T_4196 ? 16'h10 : _T_6925; // @[Mux.scala 31:69:@3823.4]
  assign _T_6927 = _T_4193 ? 16'h8 : _T_6926; // @[Mux.scala 31:69:@3824.4]
  assign _T_6928 = _T_4238 ? 16'h4 : _T_6927; // @[Mux.scala 31:69:@3825.4]
  assign _T_6929 = _T_4235 ? 16'h2 : _T_6928; // @[Mux.scala 31:69:@3826.4]
  assign _T_6930 = _T_4232 ? 16'h1 : _T_6929; // @[Mux.scala 31:69:@3827.4]
  assign _T_6931 = _T_6930[0]; // @[OneHot.scala 66:30:@3828.4]
  assign _T_6932 = _T_6930[1]; // @[OneHot.scala 66:30:@3829.4]
  assign _T_6933 = _T_6930[2]; // @[OneHot.scala 66:30:@3830.4]
  assign _T_6934 = _T_6930[3]; // @[OneHot.scala 66:30:@3831.4]
  assign _T_6935 = _T_6930[4]; // @[OneHot.scala 66:30:@3832.4]
  assign _T_6936 = _T_6930[5]; // @[OneHot.scala 66:30:@3833.4]
  assign _T_6937 = _T_6930[6]; // @[OneHot.scala 66:30:@3834.4]
  assign _T_6938 = _T_6930[7]; // @[OneHot.scala 66:30:@3835.4]
  assign _T_6939 = _T_6930[8]; // @[OneHot.scala 66:30:@3836.4]
  assign _T_6940 = _T_6930[9]; // @[OneHot.scala 66:30:@3837.4]
  assign _T_6941 = _T_6930[10]; // @[OneHot.scala 66:30:@3838.4]
  assign _T_6942 = _T_6930[11]; // @[OneHot.scala 66:30:@3839.4]
  assign _T_6943 = _T_6930[12]; // @[OneHot.scala 66:30:@3840.4]
  assign _T_6944 = _T_6930[13]; // @[OneHot.scala 66:30:@3841.4]
  assign _T_6945 = _T_6930[14]; // @[OneHot.scala 66:30:@3842.4]
  assign _T_6946 = _T_6930[15]; // @[OneHot.scala 66:30:@3843.4]
  assign _T_6987 = _T_4232 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3861.4]
  assign _T_6988 = _T_4229 ? 16'h4000 : _T_6987; // @[Mux.scala 31:69:@3862.4]
  assign _T_6989 = _T_4226 ? 16'h2000 : _T_6988; // @[Mux.scala 31:69:@3863.4]
  assign _T_6990 = _T_4223 ? 16'h1000 : _T_6989; // @[Mux.scala 31:69:@3864.4]
  assign _T_6991 = _T_4220 ? 16'h800 : _T_6990; // @[Mux.scala 31:69:@3865.4]
  assign _T_6992 = _T_4217 ? 16'h400 : _T_6991; // @[Mux.scala 31:69:@3866.4]
  assign _T_6993 = _T_4214 ? 16'h200 : _T_6992; // @[Mux.scala 31:69:@3867.4]
  assign _T_6994 = _T_4211 ? 16'h100 : _T_6993; // @[Mux.scala 31:69:@3868.4]
  assign _T_6995 = _T_4208 ? 16'h80 : _T_6994; // @[Mux.scala 31:69:@3869.4]
  assign _T_6996 = _T_4205 ? 16'h40 : _T_6995; // @[Mux.scala 31:69:@3870.4]
  assign _T_6997 = _T_4202 ? 16'h20 : _T_6996; // @[Mux.scala 31:69:@3871.4]
  assign _T_6998 = _T_4199 ? 16'h10 : _T_6997; // @[Mux.scala 31:69:@3872.4]
  assign _T_6999 = _T_4196 ? 16'h8 : _T_6998; // @[Mux.scala 31:69:@3873.4]
  assign _T_7000 = _T_4193 ? 16'h4 : _T_6999; // @[Mux.scala 31:69:@3874.4]
  assign _T_7001 = _T_4238 ? 16'h2 : _T_7000; // @[Mux.scala 31:69:@3875.4]
  assign _T_7002 = _T_4235 ? 16'h1 : _T_7001; // @[Mux.scala 31:69:@3876.4]
  assign _T_7003 = _T_7002[0]; // @[OneHot.scala 66:30:@3877.4]
  assign _T_7004 = _T_7002[1]; // @[OneHot.scala 66:30:@3878.4]
  assign _T_7005 = _T_7002[2]; // @[OneHot.scala 66:30:@3879.4]
  assign _T_7006 = _T_7002[3]; // @[OneHot.scala 66:30:@3880.4]
  assign _T_7007 = _T_7002[4]; // @[OneHot.scala 66:30:@3881.4]
  assign _T_7008 = _T_7002[5]; // @[OneHot.scala 66:30:@3882.4]
  assign _T_7009 = _T_7002[6]; // @[OneHot.scala 66:30:@3883.4]
  assign _T_7010 = _T_7002[7]; // @[OneHot.scala 66:30:@3884.4]
  assign _T_7011 = _T_7002[8]; // @[OneHot.scala 66:30:@3885.4]
  assign _T_7012 = _T_7002[9]; // @[OneHot.scala 66:30:@3886.4]
  assign _T_7013 = _T_7002[10]; // @[OneHot.scala 66:30:@3887.4]
  assign _T_7014 = _T_7002[11]; // @[OneHot.scala 66:30:@3888.4]
  assign _T_7015 = _T_7002[12]; // @[OneHot.scala 66:30:@3889.4]
  assign _T_7016 = _T_7002[13]; // @[OneHot.scala 66:30:@3890.4]
  assign _T_7017 = _T_7002[14]; // @[OneHot.scala 66:30:@3891.4]
  assign _T_7018 = _T_7002[15]; // @[OneHot.scala 66:30:@3892.4]
  assign _T_7059 = _T_4235 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3910.4]
  assign _T_7060 = _T_4232 ? 16'h4000 : _T_7059; // @[Mux.scala 31:69:@3911.4]
  assign _T_7061 = _T_4229 ? 16'h2000 : _T_7060; // @[Mux.scala 31:69:@3912.4]
  assign _T_7062 = _T_4226 ? 16'h1000 : _T_7061; // @[Mux.scala 31:69:@3913.4]
  assign _T_7063 = _T_4223 ? 16'h800 : _T_7062; // @[Mux.scala 31:69:@3914.4]
  assign _T_7064 = _T_4220 ? 16'h400 : _T_7063; // @[Mux.scala 31:69:@3915.4]
  assign _T_7065 = _T_4217 ? 16'h200 : _T_7064; // @[Mux.scala 31:69:@3916.4]
  assign _T_7066 = _T_4214 ? 16'h100 : _T_7065; // @[Mux.scala 31:69:@3917.4]
  assign _T_7067 = _T_4211 ? 16'h80 : _T_7066; // @[Mux.scala 31:69:@3918.4]
  assign _T_7068 = _T_4208 ? 16'h40 : _T_7067; // @[Mux.scala 31:69:@3919.4]
  assign _T_7069 = _T_4205 ? 16'h20 : _T_7068; // @[Mux.scala 31:69:@3920.4]
  assign _T_7070 = _T_4202 ? 16'h10 : _T_7069; // @[Mux.scala 31:69:@3921.4]
  assign _T_7071 = _T_4199 ? 16'h8 : _T_7070; // @[Mux.scala 31:69:@3922.4]
  assign _T_7072 = _T_4196 ? 16'h4 : _T_7071; // @[Mux.scala 31:69:@3923.4]
  assign _T_7073 = _T_4193 ? 16'h2 : _T_7072; // @[Mux.scala 31:69:@3924.4]
  assign _T_7074 = _T_4238 ? 16'h1 : _T_7073; // @[Mux.scala 31:69:@3925.4]
  assign _T_7075 = _T_7074[0]; // @[OneHot.scala 66:30:@3926.4]
  assign _T_7076 = _T_7074[1]; // @[OneHot.scala 66:30:@3927.4]
  assign _T_7077 = _T_7074[2]; // @[OneHot.scala 66:30:@3928.4]
  assign _T_7078 = _T_7074[3]; // @[OneHot.scala 66:30:@3929.4]
  assign _T_7079 = _T_7074[4]; // @[OneHot.scala 66:30:@3930.4]
  assign _T_7080 = _T_7074[5]; // @[OneHot.scala 66:30:@3931.4]
  assign _T_7081 = _T_7074[6]; // @[OneHot.scala 66:30:@3932.4]
  assign _T_7082 = _T_7074[7]; // @[OneHot.scala 66:30:@3933.4]
  assign _T_7083 = _T_7074[8]; // @[OneHot.scala 66:30:@3934.4]
  assign _T_7084 = _T_7074[9]; // @[OneHot.scala 66:30:@3935.4]
  assign _T_7085 = _T_7074[10]; // @[OneHot.scala 66:30:@3936.4]
  assign _T_7086 = _T_7074[11]; // @[OneHot.scala 66:30:@3937.4]
  assign _T_7087 = _T_7074[12]; // @[OneHot.scala 66:30:@3938.4]
  assign _T_7088 = _T_7074[13]; // @[OneHot.scala 66:30:@3939.4]
  assign _T_7089 = _T_7074[14]; // @[OneHot.scala 66:30:@3940.4]
  assign _T_7090 = _T_7074[15]; // @[OneHot.scala 66:30:@3941.4]
  assign _T_7155 = {_T_6002,_T_6001,_T_6000,_T_5999,_T_5998,_T_5997,_T_5996,_T_5995}; // @[Mux.scala 19:72:@3965.4]
  assign _T_7163 = {_T_6010,_T_6009,_T_6008,_T_6007,_T_6006,_T_6005,_T_6004,_T_6003,_T_7155}; // @[Mux.scala 19:72:@3973.4]
  assign _T_7165 = _T_4265 ? _T_7163 : 16'h0; // @[Mux.scala 19:72:@3974.4]
  assign _T_7172 = {_T_6073,_T_6072,_T_6071,_T_6070,_T_6069,_T_6068,_T_6067,_T_6082}; // @[Mux.scala 19:72:@3981.4]
  assign _T_7180 = {_T_6081,_T_6080,_T_6079,_T_6078,_T_6077,_T_6076,_T_6075,_T_6074,_T_7172}; // @[Mux.scala 19:72:@3989.4]
  assign _T_7182 = _T_4266 ? _T_7180 : 16'h0; // @[Mux.scala 19:72:@3990.4]
  assign _T_7189 = {_T_6144,_T_6143,_T_6142,_T_6141,_T_6140,_T_6139,_T_6154,_T_6153}; // @[Mux.scala 19:72:@3997.4]
  assign _T_7197 = {_T_6152,_T_6151,_T_6150,_T_6149,_T_6148,_T_6147,_T_6146,_T_6145,_T_7189}; // @[Mux.scala 19:72:@4005.4]
  assign _T_7199 = _T_4267 ? _T_7197 : 16'h0; // @[Mux.scala 19:72:@4006.4]
  assign _T_7206 = {_T_6215,_T_6214,_T_6213,_T_6212,_T_6211,_T_6226,_T_6225,_T_6224}; // @[Mux.scala 19:72:@4013.4]
  assign _T_7214 = {_T_6223,_T_6222,_T_6221,_T_6220,_T_6219,_T_6218,_T_6217,_T_6216,_T_7206}; // @[Mux.scala 19:72:@4021.4]
  assign _T_7216 = _T_4268 ? _T_7214 : 16'h0; // @[Mux.scala 19:72:@4022.4]
  assign _T_7223 = {_T_6286,_T_6285,_T_6284,_T_6283,_T_6298,_T_6297,_T_6296,_T_6295}; // @[Mux.scala 19:72:@4029.4]
  assign _T_7231 = {_T_6294,_T_6293,_T_6292,_T_6291,_T_6290,_T_6289,_T_6288,_T_6287,_T_7223}; // @[Mux.scala 19:72:@4037.4]
  assign _T_7233 = _T_4269 ? _T_7231 : 16'h0; // @[Mux.scala 19:72:@4038.4]
  assign _T_7240 = {_T_6357,_T_6356,_T_6355,_T_6370,_T_6369,_T_6368,_T_6367,_T_6366}; // @[Mux.scala 19:72:@4045.4]
  assign _T_7248 = {_T_6365,_T_6364,_T_6363,_T_6362,_T_6361,_T_6360,_T_6359,_T_6358,_T_7240}; // @[Mux.scala 19:72:@4053.4]
  assign _T_7250 = _T_4270 ? _T_7248 : 16'h0; // @[Mux.scala 19:72:@4054.4]
  assign _T_7257 = {_T_6428,_T_6427,_T_6442,_T_6441,_T_6440,_T_6439,_T_6438,_T_6437}; // @[Mux.scala 19:72:@4061.4]
  assign _T_7265 = {_T_6436,_T_6435,_T_6434,_T_6433,_T_6432,_T_6431,_T_6430,_T_6429,_T_7257}; // @[Mux.scala 19:72:@4069.4]
  assign _T_7267 = _T_4271 ? _T_7265 : 16'h0; // @[Mux.scala 19:72:@4070.4]
  assign _T_7274 = {_T_6499,_T_6514,_T_6513,_T_6512,_T_6511,_T_6510,_T_6509,_T_6508}; // @[Mux.scala 19:72:@4077.4]
  assign _T_7282 = {_T_6507,_T_6506,_T_6505,_T_6504,_T_6503,_T_6502,_T_6501,_T_6500,_T_7274}; // @[Mux.scala 19:72:@4085.4]
  assign _T_7284 = _T_4272 ? _T_7282 : 16'h0; // @[Mux.scala 19:72:@4086.4]
  assign _T_7291 = {_T_6586,_T_6585,_T_6584,_T_6583,_T_6582,_T_6581,_T_6580,_T_6579}; // @[Mux.scala 19:72:@4093.4]
  assign _T_7299 = {_T_6578,_T_6577,_T_6576,_T_6575,_T_6574,_T_6573,_T_6572,_T_6571,_T_7291}; // @[Mux.scala 19:72:@4101.4]
  assign _T_7301 = _T_4273 ? _T_7299 : 16'h0; // @[Mux.scala 19:72:@4102.4]
  assign _T_7308 = {_T_6657,_T_6656,_T_6655,_T_6654,_T_6653,_T_6652,_T_6651,_T_6650}; // @[Mux.scala 19:72:@4109.4]
  assign _T_7316 = {_T_6649,_T_6648,_T_6647,_T_6646,_T_6645,_T_6644,_T_6643,_T_6658,_T_7308}; // @[Mux.scala 19:72:@4117.4]
  assign _T_7318 = _T_4274 ? _T_7316 : 16'h0; // @[Mux.scala 19:72:@4118.4]
  assign _T_7325 = {_T_6728,_T_6727,_T_6726,_T_6725,_T_6724,_T_6723,_T_6722,_T_6721}; // @[Mux.scala 19:72:@4125.4]
  assign _T_7333 = {_T_6720,_T_6719,_T_6718,_T_6717,_T_6716,_T_6715,_T_6730,_T_6729,_T_7325}; // @[Mux.scala 19:72:@4133.4]
  assign _T_7335 = _T_4275 ? _T_7333 : 16'h0; // @[Mux.scala 19:72:@4134.4]
  assign _T_7342 = {_T_6799,_T_6798,_T_6797,_T_6796,_T_6795,_T_6794,_T_6793,_T_6792}; // @[Mux.scala 19:72:@4141.4]
  assign _T_7350 = {_T_6791,_T_6790,_T_6789,_T_6788,_T_6787,_T_6802,_T_6801,_T_6800,_T_7342}; // @[Mux.scala 19:72:@4149.4]
  assign _T_7352 = _T_4276 ? _T_7350 : 16'h0; // @[Mux.scala 19:72:@4150.4]
  assign _T_7359 = {_T_6870,_T_6869,_T_6868,_T_6867,_T_6866,_T_6865,_T_6864,_T_6863}; // @[Mux.scala 19:72:@4157.4]
  assign _T_7367 = {_T_6862,_T_6861,_T_6860,_T_6859,_T_6874,_T_6873,_T_6872,_T_6871,_T_7359}; // @[Mux.scala 19:72:@4165.4]
  assign _T_7369 = _T_4277 ? _T_7367 : 16'h0; // @[Mux.scala 19:72:@4166.4]
  assign _T_7376 = {_T_6941,_T_6940,_T_6939,_T_6938,_T_6937,_T_6936,_T_6935,_T_6934}; // @[Mux.scala 19:72:@4173.4]
  assign _T_7384 = {_T_6933,_T_6932,_T_6931,_T_6946,_T_6945,_T_6944,_T_6943,_T_6942,_T_7376}; // @[Mux.scala 19:72:@4181.4]
  assign _T_7386 = _T_4278 ? _T_7384 : 16'h0; // @[Mux.scala 19:72:@4182.4]
  assign _T_7393 = {_T_7012,_T_7011,_T_7010,_T_7009,_T_7008,_T_7007,_T_7006,_T_7005}; // @[Mux.scala 19:72:@4189.4]
  assign _T_7401 = {_T_7004,_T_7003,_T_7018,_T_7017,_T_7016,_T_7015,_T_7014,_T_7013,_T_7393}; // @[Mux.scala 19:72:@4197.4]
  assign _T_7403 = _T_4279 ? _T_7401 : 16'h0; // @[Mux.scala 19:72:@4198.4]
  assign _T_7410 = {_T_7083,_T_7082,_T_7081,_T_7080,_T_7079,_T_7078,_T_7077,_T_7076}; // @[Mux.scala 19:72:@4205.4]
  assign _T_7418 = {_T_7075,_T_7090,_T_7089,_T_7088,_T_7087,_T_7086,_T_7085,_T_7084,_T_7410}; // @[Mux.scala 19:72:@4213.4]
  assign _T_7420 = _T_4280 ? _T_7418 : 16'h0; // @[Mux.scala 19:72:@4214.4]
  assign _T_7421 = _T_7165 | _T_7182; // @[Mux.scala 19:72:@4215.4]
  assign _T_7422 = _T_7421 | _T_7199; // @[Mux.scala 19:72:@4216.4]
  assign _T_7423 = _T_7422 | _T_7216; // @[Mux.scala 19:72:@4217.4]
  assign _T_7424 = _T_7423 | _T_7233; // @[Mux.scala 19:72:@4218.4]
  assign _T_7425 = _T_7424 | _T_7250; // @[Mux.scala 19:72:@4219.4]
  assign _T_7426 = _T_7425 | _T_7267; // @[Mux.scala 19:72:@4220.4]
  assign _T_7427 = _T_7426 | _T_7284; // @[Mux.scala 19:72:@4221.4]
  assign _T_7428 = _T_7427 | _T_7301; // @[Mux.scala 19:72:@4222.4]
  assign _T_7429 = _T_7428 | _T_7318; // @[Mux.scala 19:72:@4223.4]
  assign _T_7430 = _T_7429 | _T_7335; // @[Mux.scala 19:72:@4224.4]
  assign _T_7431 = _T_7430 | _T_7352; // @[Mux.scala 19:72:@4225.4]
  assign _T_7432 = _T_7431 | _T_7369; // @[Mux.scala 19:72:@4226.4]
  assign _T_7433 = _T_7432 | _T_7386; // @[Mux.scala 19:72:@4227.4]
  assign _T_7434 = _T_7433 | _T_7403; // @[Mux.scala 19:72:@4228.4]
  assign _T_7435 = _T_7434 | _T_7420; // @[Mux.scala 19:72:@4229.4]
  assign inputDataPriorityPorts_0_0 = _T_7435[0]; // @[Mux.scala 19:72:@4233.4]
  assign inputDataPriorityPorts_0_1 = _T_7435[1]; // @[Mux.scala 19:72:@4235.4]
  assign inputDataPriorityPorts_0_2 = _T_7435[2]; // @[Mux.scala 19:72:@4237.4]
  assign inputDataPriorityPorts_0_3 = _T_7435[3]; // @[Mux.scala 19:72:@4239.4]
  assign inputDataPriorityPorts_0_4 = _T_7435[4]; // @[Mux.scala 19:72:@4241.4]
  assign inputDataPriorityPorts_0_5 = _T_7435[5]; // @[Mux.scala 19:72:@4243.4]
  assign inputDataPriorityPorts_0_6 = _T_7435[6]; // @[Mux.scala 19:72:@4245.4]
  assign inputDataPriorityPorts_0_7 = _T_7435[7]; // @[Mux.scala 19:72:@4247.4]
  assign inputDataPriorityPorts_0_8 = _T_7435[8]; // @[Mux.scala 19:72:@4249.4]
  assign inputDataPriorityPorts_0_9 = _T_7435[9]; // @[Mux.scala 19:72:@4251.4]
  assign inputDataPriorityPorts_0_10 = _T_7435[10]; // @[Mux.scala 19:72:@4253.4]
  assign inputDataPriorityPorts_0_11 = _T_7435[11]; // @[Mux.scala 19:72:@4255.4]
  assign inputDataPriorityPorts_0_12 = _T_7435[12]; // @[Mux.scala 19:72:@4257.4]
  assign inputDataPriorityPorts_0_13 = _T_7435[13]; // @[Mux.scala 19:72:@4259.4]
  assign inputDataPriorityPorts_0_14 = _T_7435[14]; // @[Mux.scala 19:72:@4261.4]
  assign inputDataPriorityPorts_0_15 = _T_7435[15]; // @[Mux.scala 19:72:@4263.4]
  assign _T_7581 = inputAddrPriorityPorts_0_0 & _T_4122; // @[StoreQueue.scala 209:52:@4287.6]
  assign _T_7582 = _T_7581 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4288.6]
  assign _GEN_992 = _T_7582 ? io_addressFromStorePorts_0 : addrQ_0; // @[StoreQueue.scala 210:40:@4292.6]
  assign _GEN_993 = _T_7582 ? 1'h1 : addrKnown_0; // @[StoreQueue.scala 210:40:@4292.6]
  assign _T_7598 = inputDataPriorityPorts_0_0 & _T_4192; // @[StoreQueue.scala 215:52:@4297.6]
  assign _T_7599 = _T_7598 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4298.6]
  assign _GEN_994 = _T_7599 ? io_dataFromStorePorts_0 : dataQ_0; // @[StoreQueue.scala 216:40:@4302.6]
  assign _GEN_995 = _T_7599 ? 1'h1 : dataKnown_0; // @[StoreQueue.scala 216:40:@4302.6]
  assign _GEN_996 = initBits_0 ? 1'h0 : _GEN_993; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_997 = initBits_0 ? 1'h0 : _GEN_995; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_998 = initBits_0 ? addrQ_0 : _GEN_992; // @[StoreQueue.scala 204:35:@4281.4]
  assign _GEN_999 = initBits_0 ? dataQ_0 : _GEN_994; // @[StoreQueue.scala 204:35:@4281.4]
  assign _T_7617 = inputAddrPriorityPorts_0_1 & _T_4125; // @[StoreQueue.scala 209:52:@4313.6]
  assign _T_7618 = _T_7617 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4314.6]
  assign _GEN_1000 = _T_7618 ? io_addressFromStorePorts_0 : addrQ_1; // @[StoreQueue.scala 210:40:@4318.6]
  assign _GEN_1001 = _T_7618 ? 1'h1 : addrKnown_1; // @[StoreQueue.scala 210:40:@4318.6]
  assign _T_7634 = inputDataPriorityPorts_0_1 & _T_4195; // @[StoreQueue.scala 215:52:@4323.6]
  assign _T_7635 = _T_7634 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4324.6]
  assign _GEN_1002 = _T_7635 ? io_dataFromStorePorts_0 : dataQ_1; // @[StoreQueue.scala 216:40:@4328.6]
  assign _GEN_1003 = _T_7635 ? 1'h1 : dataKnown_1; // @[StoreQueue.scala 216:40:@4328.6]
  assign _GEN_1004 = initBits_1 ? 1'h0 : _GEN_1001; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1005 = initBits_1 ? 1'h0 : _GEN_1003; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1006 = initBits_1 ? addrQ_1 : _GEN_1000; // @[StoreQueue.scala 204:35:@4307.4]
  assign _GEN_1007 = initBits_1 ? dataQ_1 : _GEN_1002; // @[StoreQueue.scala 204:35:@4307.4]
  assign _T_7653 = inputAddrPriorityPorts_0_2 & _T_4128; // @[StoreQueue.scala 209:52:@4339.6]
  assign _T_7654 = _T_7653 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4340.6]
  assign _GEN_1008 = _T_7654 ? io_addressFromStorePorts_0 : addrQ_2; // @[StoreQueue.scala 210:40:@4344.6]
  assign _GEN_1009 = _T_7654 ? 1'h1 : addrKnown_2; // @[StoreQueue.scala 210:40:@4344.6]
  assign _T_7670 = inputDataPriorityPorts_0_2 & _T_4198; // @[StoreQueue.scala 215:52:@4349.6]
  assign _T_7671 = _T_7670 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4350.6]
  assign _GEN_1010 = _T_7671 ? io_dataFromStorePorts_0 : dataQ_2; // @[StoreQueue.scala 216:40:@4354.6]
  assign _GEN_1011 = _T_7671 ? 1'h1 : dataKnown_2; // @[StoreQueue.scala 216:40:@4354.6]
  assign _GEN_1012 = initBits_2 ? 1'h0 : _GEN_1009; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1013 = initBits_2 ? 1'h0 : _GEN_1011; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1014 = initBits_2 ? addrQ_2 : _GEN_1008; // @[StoreQueue.scala 204:35:@4333.4]
  assign _GEN_1015 = initBits_2 ? dataQ_2 : _GEN_1010; // @[StoreQueue.scala 204:35:@4333.4]
  assign _T_7689 = inputAddrPriorityPorts_0_3 & _T_4131; // @[StoreQueue.scala 209:52:@4365.6]
  assign _T_7690 = _T_7689 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4366.6]
  assign _GEN_1016 = _T_7690 ? io_addressFromStorePorts_0 : addrQ_3; // @[StoreQueue.scala 210:40:@4370.6]
  assign _GEN_1017 = _T_7690 ? 1'h1 : addrKnown_3; // @[StoreQueue.scala 210:40:@4370.6]
  assign _T_7706 = inputDataPriorityPorts_0_3 & _T_4201; // @[StoreQueue.scala 215:52:@4375.6]
  assign _T_7707 = _T_7706 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4376.6]
  assign _GEN_1018 = _T_7707 ? io_dataFromStorePorts_0 : dataQ_3; // @[StoreQueue.scala 216:40:@4380.6]
  assign _GEN_1019 = _T_7707 ? 1'h1 : dataKnown_3; // @[StoreQueue.scala 216:40:@4380.6]
  assign _GEN_1020 = initBits_3 ? 1'h0 : _GEN_1017; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1021 = initBits_3 ? 1'h0 : _GEN_1019; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1022 = initBits_3 ? addrQ_3 : _GEN_1016; // @[StoreQueue.scala 204:35:@4359.4]
  assign _GEN_1023 = initBits_3 ? dataQ_3 : _GEN_1018; // @[StoreQueue.scala 204:35:@4359.4]
  assign _T_7725 = inputAddrPriorityPorts_0_4 & _T_4134; // @[StoreQueue.scala 209:52:@4391.6]
  assign _T_7726 = _T_7725 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4392.6]
  assign _GEN_1024 = _T_7726 ? io_addressFromStorePorts_0 : addrQ_4; // @[StoreQueue.scala 210:40:@4396.6]
  assign _GEN_1025 = _T_7726 ? 1'h1 : addrKnown_4; // @[StoreQueue.scala 210:40:@4396.6]
  assign _T_7742 = inputDataPriorityPorts_0_4 & _T_4204; // @[StoreQueue.scala 215:52:@4401.6]
  assign _T_7743 = _T_7742 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4402.6]
  assign _GEN_1026 = _T_7743 ? io_dataFromStorePorts_0 : dataQ_4; // @[StoreQueue.scala 216:40:@4406.6]
  assign _GEN_1027 = _T_7743 ? 1'h1 : dataKnown_4; // @[StoreQueue.scala 216:40:@4406.6]
  assign _GEN_1028 = initBits_4 ? 1'h0 : _GEN_1025; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1029 = initBits_4 ? 1'h0 : _GEN_1027; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1030 = initBits_4 ? addrQ_4 : _GEN_1024; // @[StoreQueue.scala 204:35:@4385.4]
  assign _GEN_1031 = initBits_4 ? dataQ_4 : _GEN_1026; // @[StoreQueue.scala 204:35:@4385.4]
  assign _T_7761 = inputAddrPriorityPorts_0_5 & _T_4137; // @[StoreQueue.scala 209:52:@4417.6]
  assign _T_7762 = _T_7761 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4418.6]
  assign _GEN_1032 = _T_7762 ? io_addressFromStorePorts_0 : addrQ_5; // @[StoreQueue.scala 210:40:@4422.6]
  assign _GEN_1033 = _T_7762 ? 1'h1 : addrKnown_5; // @[StoreQueue.scala 210:40:@4422.6]
  assign _T_7778 = inputDataPriorityPorts_0_5 & _T_4207; // @[StoreQueue.scala 215:52:@4427.6]
  assign _T_7779 = _T_7778 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4428.6]
  assign _GEN_1034 = _T_7779 ? io_dataFromStorePorts_0 : dataQ_5; // @[StoreQueue.scala 216:40:@4432.6]
  assign _GEN_1035 = _T_7779 ? 1'h1 : dataKnown_5; // @[StoreQueue.scala 216:40:@4432.6]
  assign _GEN_1036 = initBits_5 ? 1'h0 : _GEN_1033; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1037 = initBits_5 ? 1'h0 : _GEN_1035; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1038 = initBits_5 ? addrQ_5 : _GEN_1032; // @[StoreQueue.scala 204:35:@4411.4]
  assign _GEN_1039 = initBits_5 ? dataQ_5 : _GEN_1034; // @[StoreQueue.scala 204:35:@4411.4]
  assign _T_7797 = inputAddrPriorityPorts_0_6 & _T_4140; // @[StoreQueue.scala 209:52:@4443.6]
  assign _T_7798 = _T_7797 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4444.6]
  assign _GEN_1040 = _T_7798 ? io_addressFromStorePorts_0 : addrQ_6; // @[StoreQueue.scala 210:40:@4448.6]
  assign _GEN_1041 = _T_7798 ? 1'h1 : addrKnown_6; // @[StoreQueue.scala 210:40:@4448.6]
  assign _T_7814 = inputDataPriorityPorts_0_6 & _T_4210; // @[StoreQueue.scala 215:52:@4453.6]
  assign _T_7815 = _T_7814 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4454.6]
  assign _GEN_1042 = _T_7815 ? io_dataFromStorePorts_0 : dataQ_6; // @[StoreQueue.scala 216:40:@4458.6]
  assign _GEN_1043 = _T_7815 ? 1'h1 : dataKnown_6; // @[StoreQueue.scala 216:40:@4458.6]
  assign _GEN_1044 = initBits_6 ? 1'h0 : _GEN_1041; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1045 = initBits_6 ? 1'h0 : _GEN_1043; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1046 = initBits_6 ? addrQ_6 : _GEN_1040; // @[StoreQueue.scala 204:35:@4437.4]
  assign _GEN_1047 = initBits_6 ? dataQ_6 : _GEN_1042; // @[StoreQueue.scala 204:35:@4437.4]
  assign _T_7833 = inputAddrPriorityPorts_0_7 & _T_4143; // @[StoreQueue.scala 209:52:@4469.6]
  assign _T_7834 = _T_7833 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4470.6]
  assign _GEN_1048 = _T_7834 ? io_addressFromStorePorts_0 : addrQ_7; // @[StoreQueue.scala 210:40:@4474.6]
  assign _GEN_1049 = _T_7834 ? 1'h1 : addrKnown_7; // @[StoreQueue.scala 210:40:@4474.6]
  assign _T_7850 = inputDataPriorityPorts_0_7 & _T_4213; // @[StoreQueue.scala 215:52:@4479.6]
  assign _T_7851 = _T_7850 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4480.6]
  assign _GEN_1050 = _T_7851 ? io_dataFromStorePorts_0 : dataQ_7; // @[StoreQueue.scala 216:40:@4484.6]
  assign _GEN_1051 = _T_7851 ? 1'h1 : dataKnown_7; // @[StoreQueue.scala 216:40:@4484.6]
  assign _GEN_1052 = initBits_7 ? 1'h0 : _GEN_1049; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1053 = initBits_7 ? 1'h0 : _GEN_1051; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1054 = initBits_7 ? addrQ_7 : _GEN_1048; // @[StoreQueue.scala 204:35:@4463.4]
  assign _GEN_1055 = initBits_7 ? dataQ_7 : _GEN_1050; // @[StoreQueue.scala 204:35:@4463.4]
  assign _T_7869 = inputAddrPriorityPorts_0_8 & _T_4146; // @[StoreQueue.scala 209:52:@4495.6]
  assign _T_7870 = _T_7869 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4496.6]
  assign _GEN_1056 = _T_7870 ? io_addressFromStorePorts_0 : addrQ_8; // @[StoreQueue.scala 210:40:@4500.6]
  assign _GEN_1057 = _T_7870 ? 1'h1 : addrKnown_8; // @[StoreQueue.scala 210:40:@4500.6]
  assign _T_7886 = inputDataPriorityPorts_0_8 & _T_4216; // @[StoreQueue.scala 215:52:@4505.6]
  assign _T_7887 = _T_7886 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4506.6]
  assign _GEN_1058 = _T_7887 ? io_dataFromStorePorts_0 : dataQ_8; // @[StoreQueue.scala 216:40:@4510.6]
  assign _GEN_1059 = _T_7887 ? 1'h1 : dataKnown_8; // @[StoreQueue.scala 216:40:@4510.6]
  assign _GEN_1060 = initBits_8 ? 1'h0 : _GEN_1057; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1061 = initBits_8 ? 1'h0 : _GEN_1059; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1062 = initBits_8 ? addrQ_8 : _GEN_1056; // @[StoreQueue.scala 204:35:@4489.4]
  assign _GEN_1063 = initBits_8 ? dataQ_8 : _GEN_1058; // @[StoreQueue.scala 204:35:@4489.4]
  assign _T_7905 = inputAddrPriorityPorts_0_9 & _T_4149; // @[StoreQueue.scala 209:52:@4521.6]
  assign _T_7906 = _T_7905 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4522.6]
  assign _GEN_1064 = _T_7906 ? io_addressFromStorePorts_0 : addrQ_9; // @[StoreQueue.scala 210:40:@4526.6]
  assign _GEN_1065 = _T_7906 ? 1'h1 : addrKnown_9; // @[StoreQueue.scala 210:40:@4526.6]
  assign _T_7922 = inputDataPriorityPorts_0_9 & _T_4219; // @[StoreQueue.scala 215:52:@4531.6]
  assign _T_7923 = _T_7922 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4532.6]
  assign _GEN_1066 = _T_7923 ? io_dataFromStorePorts_0 : dataQ_9; // @[StoreQueue.scala 216:40:@4536.6]
  assign _GEN_1067 = _T_7923 ? 1'h1 : dataKnown_9; // @[StoreQueue.scala 216:40:@4536.6]
  assign _GEN_1068 = initBits_9 ? 1'h0 : _GEN_1065; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1069 = initBits_9 ? 1'h0 : _GEN_1067; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1070 = initBits_9 ? addrQ_9 : _GEN_1064; // @[StoreQueue.scala 204:35:@4515.4]
  assign _GEN_1071 = initBits_9 ? dataQ_9 : _GEN_1066; // @[StoreQueue.scala 204:35:@4515.4]
  assign _T_7941 = inputAddrPriorityPorts_0_10 & _T_4152; // @[StoreQueue.scala 209:52:@4547.6]
  assign _T_7942 = _T_7941 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4548.6]
  assign _GEN_1072 = _T_7942 ? io_addressFromStorePorts_0 : addrQ_10; // @[StoreQueue.scala 210:40:@4552.6]
  assign _GEN_1073 = _T_7942 ? 1'h1 : addrKnown_10; // @[StoreQueue.scala 210:40:@4552.6]
  assign _T_7958 = inputDataPriorityPorts_0_10 & _T_4222; // @[StoreQueue.scala 215:52:@4557.6]
  assign _T_7959 = _T_7958 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4558.6]
  assign _GEN_1074 = _T_7959 ? io_dataFromStorePorts_0 : dataQ_10; // @[StoreQueue.scala 216:40:@4562.6]
  assign _GEN_1075 = _T_7959 ? 1'h1 : dataKnown_10; // @[StoreQueue.scala 216:40:@4562.6]
  assign _GEN_1076 = initBits_10 ? 1'h0 : _GEN_1073; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1077 = initBits_10 ? 1'h0 : _GEN_1075; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1078 = initBits_10 ? addrQ_10 : _GEN_1072; // @[StoreQueue.scala 204:35:@4541.4]
  assign _GEN_1079 = initBits_10 ? dataQ_10 : _GEN_1074; // @[StoreQueue.scala 204:35:@4541.4]
  assign _T_7977 = inputAddrPriorityPorts_0_11 & _T_4155; // @[StoreQueue.scala 209:52:@4573.6]
  assign _T_7978 = _T_7977 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4574.6]
  assign _GEN_1080 = _T_7978 ? io_addressFromStorePorts_0 : addrQ_11; // @[StoreQueue.scala 210:40:@4578.6]
  assign _GEN_1081 = _T_7978 ? 1'h1 : addrKnown_11; // @[StoreQueue.scala 210:40:@4578.6]
  assign _T_7994 = inputDataPriorityPorts_0_11 & _T_4225; // @[StoreQueue.scala 215:52:@4583.6]
  assign _T_7995 = _T_7994 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4584.6]
  assign _GEN_1082 = _T_7995 ? io_dataFromStorePorts_0 : dataQ_11; // @[StoreQueue.scala 216:40:@4588.6]
  assign _GEN_1083 = _T_7995 ? 1'h1 : dataKnown_11; // @[StoreQueue.scala 216:40:@4588.6]
  assign _GEN_1084 = initBits_11 ? 1'h0 : _GEN_1081; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1085 = initBits_11 ? 1'h0 : _GEN_1083; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1086 = initBits_11 ? addrQ_11 : _GEN_1080; // @[StoreQueue.scala 204:35:@4567.4]
  assign _GEN_1087 = initBits_11 ? dataQ_11 : _GEN_1082; // @[StoreQueue.scala 204:35:@4567.4]
  assign _T_8013 = inputAddrPriorityPorts_0_12 & _T_4158; // @[StoreQueue.scala 209:52:@4599.6]
  assign _T_8014 = _T_8013 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4600.6]
  assign _GEN_1088 = _T_8014 ? io_addressFromStorePorts_0 : addrQ_12; // @[StoreQueue.scala 210:40:@4604.6]
  assign _GEN_1089 = _T_8014 ? 1'h1 : addrKnown_12; // @[StoreQueue.scala 210:40:@4604.6]
  assign _T_8030 = inputDataPriorityPorts_0_12 & _T_4228; // @[StoreQueue.scala 215:52:@4609.6]
  assign _T_8031 = _T_8030 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4610.6]
  assign _GEN_1090 = _T_8031 ? io_dataFromStorePorts_0 : dataQ_12; // @[StoreQueue.scala 216:40:@4614.6]
  assign _GEN_1091 = _T_8031 ? 1'h1 : dataKnown_12; // @[StoreQueue.scala 216:40:@4614.6]
  assign _GEN_1092 = initBits_12 ? 1'h0 : _GEN_1089; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1093 = initBits_12 ? 1'h0 : _GEN_1091; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1094 = initBits_12 ? addrQ_12 : _GEN_1088; // @[StoreQueue.scala 204:35:@4593.4]
  assign _GEN_1095 = initBits_12 ? dataQ_12 : _GEN_1090; // @[StoreQueue.scala 204:35:@4593.4]
  assign _T_8049 = inputAddrPriorityPorts_0_13 & _T_4161; // @[StoreQueue.scala 209:52:@4625.6]
  assign _T_8050 = _T_8049 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4626.6]
  assign _GEN_1096 = _T_8050 ? io_addressFromStorePorts_0 : addrQ_13; // @[StoreQueue.scala 210:40:@4630.6]
  assign _GEN_1097 = _T_8050 ? 1'h1 : addrKnown_13; // @[StoreQueue.scala 210:40:@4630.6]
  assign _T_8066 = inputDataPriorityPorts_0_13 & _T_4231; // @[StoreQueue.scala 215:52:@4635.6]
  assign _T_8067 = _T_8066 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4636.6]
  assign _GEN_1098 = _T_8067 ? io_dataFromStorePorts_0 : dataQ_13; // @[StoreQueue.scala 216:40:@4640.6]
  assign _GEN_1099 = _T_8067 ? 1'h1 : dataKnown_13; // @[StoreQueue.scala 216:40:@4640.6]
  assign _GEN_1100 = initBits_13 ? 1'h0 : _GEN_1097; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1101 = initBits_13 ? 1'h0 : _GEN_1099; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1102 = initBits_13 ? addrQ_13 : _GEN_1096; // @[StoreQueue.scala 204:35:@4619.4]
  assign _GEN_1103 = initBits_13 ? dataQ_13 : _GEN_1098; // @[StoreQueue.scala 204:35:@4619.4]
  assign _T_8085 = inputAddrPriorityPorts_0_14 & _T_4164; // @[StoreQueue.scala 209:52:@4651.6]
  assign _T_8086 = _T_8085 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4652.6]
  assign _GEN_1104 = _T_8086 ? io_addressFromStorePorts_0 : addrQ_14; // @[StoreQueue.scala 210:40:@4656.6]
  assign _GEN_1105 = _T_8086 ? 1'h1 : addrKnown_14; // @[StoreQueue.scala 210:40:@4656.6]
  assign _T_8102 = inputDataPriorityPorts_0_14 & _T_4234; // @[StoreQueue.scala 215:52:@4661.6]
  assign _T_8103 = _T_8102 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4662.6]
  assign _GEN_1106 = _T_8103 ? io_dataFromStorePorts_0 : dataQ_14; // @[StoreQueue.scala 216:40:@4666.6]
  assign _GEN_1107 = _T_8103 ? 1'h1 : dataKnown_14; // @[StoreQueue.scala 216:40:@4666.6]
  assign _GEN_1108 = initBits_14 ? 1'h0 : _GEN_1105; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1109 = initBits_14 ? 1'h0 : _GEN_1107; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1110 = initBits_14 ? addrQ_14 : _GEN_1104; // @[StoreQueue.scala 204:35:@4645.4]
  assign _GEN_1111 = initBits_14 ? dataQ_14 : _GEN_1106; // @[StoreQueue.scala 204:35:@4645.4]
  assign _T_8121 = inputAddrPriorityPorts_0_15 & _T_4167; // @[StoreQueue.scala 209:52:@4677.6]
  assign _T_8122 = _T_8121 & io_storeAddrEnable_0; // @[StoreQueue.scala 209:81:@4678.6]
  assign _GEN_1112 = _T_8122 ? io_addressFromStorePorts_0 : addrQ_15; // @[StoreQueue.scala 210:40:@4682.6]
  assign _GEN_1113 = _T_8122 ? 1'h1 : addrKnown_15; // @[StoreQueue.scala 210:40:@4682.6]
  assign _T_8138 = inputDataPriorityPorts_0_15 & _T_4237; // @[StoreQueue.scala 215:52:@4687.6]
  assign _T_8139 = _T_8138 & io_storeDataEnable_0; // @[StoreQueue.scala 215:81:@4688.6]
  assign _GEN_1114 = _T_8139 ? io_dataFromStorePorts_0 : dataQ_15; // @[StoreQueue.scala 216:40:@4692.6]
  assign _GEN_1115 = _T_8139 ? 1'h1 : dataKnown_15; // @[StoreQueue.scala 216:40:@4692.6]
  assign _GEN_1116 = initBits_15 ? 1'h0 : _GEN_1113; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1117 = initBits_15 ? 1'h0 : _GEN_1115; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1118 = initBits_15 ? addrQ_15 : _GEN_1112; // @[StoreQueue.scala 204:35:@4671.4]
  assign _GEN_1119 = initBits_15 ? dataQ_15 : _GEN_1114; // @[StoreQueue.scala 204:35:@4671.4]
  assign _T_8153 = storeRequest & io_memIsReadyForStores; // @[StoreQueue.scala 229:23:@4697.4]
  assign _T_8156 = head + 4'h1; // @[util.scala 10:8:@4699.6]
  assign _GEN_64 = _T_8156 % 5'h10; // @[util.scala 10:14:@4700.6]
  assign _T_8157 = _GEN_64[4:0]; // @[util.scala 10:14:@4700.6]
  assign _GEN_1120 = _T_8153 ? _T_8157 : {{1'd0}, head}; // @[StoreQueue.scala 229:50:@4698.4]
  assign _GEN_1234 = {{3'd0}, io_bbNumStores}; // @[util.scala 10:8:@4704.6]
  assign _T_8159 = tail + _GEN_1234; // @[util.scala 10:8:@4704.6]
  assign _GEN_65 = _T_8159 % 5'h10; // @[util.scala 10:14:@4705.6]
  assign _T_8160 = _GEN_65[4:0]; // @[util.scala 10:14:@4705.6]
  assign _GEN_1121 = io_bbStart ? _T_8160 : {{1'd0}, tail}; // @[StoreQueue.scala 233:20:@4703.4]
  assign _T_8162 = allocatedEntries_0 == 1'h0; // @[StoreQueue.scala 237:84:@4708.4]
  assign _T_8163 = storeCompleted_0 | _T_8162; // @[StoreQueue.scala 237:81:@4709.4]
  assign _T_8165 = allocatedEntries_1 == 1'h0; // @[StoreQueue.scala 237:84:@4710.4]
  assign _T_8166 = storeCompleted_1 | _T_8165; // @[StoreQueue.scala 237:81:@4711.4]
  assign _T_8168 = allocatedEntries_2 == 1'h0; // @[StoreQueue.scala 237:84:@4712.4]
  assign _T_8169 = storeCompleted_2 | _T_8168; // @[StoreQueue.scala 237:81:@4713.4]
  assign _T_8171 = allocatedEntries_3 == 1'h0; // @[StoreQueue.scala 237:84:@4714.4]
  assign _T_8172 = storeCompleted_3 | _T_8171; // @[StoreQueue.scala 237:81:@4715.4]
  assign _T_8174 = allocatedEntries_4 == 1'h0; // @[StoreQueue.scala 237:84:@4716.4]
  assign _T_8175 = storeCompleted_4 | _T_8174; // @[StoreQueue.scala 237:81:@4717.4]
  assign _T_8177 = allocatedEntries_5 == 1'h0; // @[StoreQueue.scala 237:84:@4718.4]
  assign _T_8178 = storeCompleted_5 | _T_8177; // @[StoreQueue.scala 237:81:@4719.4]
  assign _T_8180 = allocatedEntries_6 == 1'h0; // @[StoreQueue.scala 237:84:@4720.4]
  assign _T_8181 = storeCompleted_6 | _T_8180; // @[StoreQueue.scala 237:81:@4721.4]
  assign _T_8183 = allocatedEntries_7 == 1'h0; // @[StoreQueue.scala 237:84:@4722.4]
  assign _T_8184 = storeCompleted_7 | _T_8183; // @[StoreQueue.scala 237:81:@4723.4]
  assign _T_8186 = allocatedEntries_8 == 1'h0; // @[StoreQueue.scala 237:84:@4724.4]
  assign _T_8187 = storeCompleted_8 | _T_8186; // @[StoreQueue.scala 237:81:@4725.4]
  assign _T_8189 = allocatedEntries_9 == 1'h0; // @[StoreQueue.scala 237:84:@4726.4]
  assign _T_8190 = storeCompleted_9 | _T_8189; // @[StoreQueue.scala 237:81:@4727.4]
  assign _T_8192 = allocatedEntries_10 == 1'h0; // @[StoreQueue.scala 237:84:@4728.4]
  assign _T_8193 = storeCompleted_10 | _T_8192; // @[StoreQueue.scala 237:81:@4729.4]
  assign _T_8195 = allocatedEntries_11 == 1'h0; // @[StoreQueue.scala 237:84:@4730.4]
  assign _T_8196 = storeCompleted_11 | _T_8195; // @[StoreQueue.scala 237:81:@4731.4]
  assign _T_8198 = allocatedEntries_12 == 1'h0; // @[StoreQueue.scala 237:84:@4732.4]
  assign _T_8199 = storeCompleted_12 | _T_8198; // @[StoreQueue.scala 237:81:@4733.4]
  assign _T_8201 = allocatedEntries_13 == 1'h0; // @[StoreQueue.scala 237:84:@4734.4]
  assign _T_8202 = storeCompleted_13 | _T_8201; // @[StoreQueue.scala 237:81:@4735.4]
  assign _T_8204 = allocatedEntries_14 == 1'h0; // @[StoreQueue.scala 237:84:@4736.4]
  assign _T_8205 = storeCompleted_14 | _T_8204; // @[StoreQueue.scala 237:81:@4737.4]
  assign _T_8207 = allocatedEntries_15 == 1'h0; // @[StoreQueue.scala 237:84:@4738.4]
  assign _T_8208 = storeCompleted_15 | _T_8207; // @[StoreQueue.scala 237:81:@4739.4]
  assign _T_8233 = _T_8163 & _T_8166; // @[StoreQueue.scala 237:98:@4758.4]
  assign _T_8234 = _T_8233 & _T_8169; // @[StoreQueue.scala 237:98:@4759.4]
  assign _T_8235 = _T_8234 & _T_8172; // @[StoreQueue.scala 237:98:@4760.4]
  assign _T_8236 = _T_8235 & _T_8175; // @[StoreQueue.scala 237:98:@4761.4]
  assign _T_8237 = _T_8236 & _T_8178; // @[StoreQueue.scala 237:98:@4762.4]
  assign _T_8238 = _T_8237 & _T_8181; // @[StoreQueue.scala 237:98:@4763.4]
  assign _T_8239 = _T_8238 & _T_8184; // @[StoreQueue.scala 237:98:@4764.4]
  assign _T_8240 = _T_8239 & _T_8187; // @[StoreQueue.scala 237:98:@4765.4]
  assign _T_8241 = _T_8240 & _T_8190; // @[StoreQueue.scala 237:98:@4766.4]
  assign _T_8242 = _T_8241 & _T_8193; // @[StoreQueue.scala 237:98:@4767.4]
  assign _T_8243 = _T_8242 & _T_8196; // @[StoreQueue.scala 237:98:@4768.4]
  assign _T_8244 = _T_8243 & _T_8199; // @[StoreQueue.scala 237:98:@4769.4]
  assign _T_8245 = _T_8244 & _T_8202; // @[StoreQueue.scala 237:98:@4770.4]
  assign _T_8246 = _T_8245 & _T_8205; // @[StoreQueue.scala 237:98:@4771.4]
  assign _GEN_1123 = 4'h1 == head ? dataQ_1 : dataQ_0; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1124 = 4'h2 == head ? dataQ_2 : _GEN_1123; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1125 = 4'h3 == head ? dataQ_3 : _GEN_1124; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1126 = 4'h4 == head ? dataQ_4 : _GEN_1125; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1127 = 4'h5 == head ? dataQ_5 : _GEN_1126; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1128 = 4'h6 == head ? dataQ_6 : _GEN_1127; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1129 = 4'h7 == head ? dataQ_7 : _GEN_1128; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1130 = 4'h8 == head ? dataQ_8 : _GEN_1129; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1131 = 4'h9 == head ? dataQ_9 : _GEN_1130; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1132 = 4'ha == head ? dataQ_10 : _GEN_1131; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1133 = 4'hb == head ? dataQ_11 : _GEN_1132; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1134 = 4'hc == head ? dataQ_12 : _GEN_1133; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1135 = 4'hd == head ? dataQ_13 : _GEN_1134; // @[StoreQueue.scala 252:21:@4841.4]
  assign _GEN_1136 = 4'he == head ? dataQ_14 : _GEN_1135; // @[StoreQueue.scala 252:21:@4841.4]
  assign io_storeTail = tail; // @[StoreQueue.scala 246:16:@4775.4]
  assign io_storeHead = head; // @[StoreQueue.scala 245:16:@4774.4]
  assign io_storeEmpty = _T_8246 & _T_8208; // @[StoreQueue.scala 237:17:@4773.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[StoreQueue.scala 250:20:@4824.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[StoreQueue.scala 250:20:@4825.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[StoreQueue.scala 250:20:@4826.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[StoreQueue.scala 250:20:@4827.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[StoreQueue.scala 250:20:@4828.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[StoreQueue.scala 250:20:@4829.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[StoreQueue.scala 250:20:@4830.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[StoreQueue.scala 250:20:@4831.4]
  assign io_storeAddrDone_8 = addrKnown_8; // @[StoreQueue.scala 250:20:@4832.4]
  assign io_storeAddrDone_9 = addrKnown_9; // @[StoreQueue.scala 250:20:@4833.4]
  assign io_storeAddrDone_10 = addrKnown_10; // @[StoreQueue.scala 250:20:@4834.4]
  assign io_storeAddrDone_11 = addrKnown_11; // @[StoreQueue.scala 250:20:@4835.4]
  assign io_storeAddrDone_12 = addrKnown_12; // @[StoreQueue.scala 250:20:@4836.4]
  assign io_storeAddrDone_13 = addrKnown_13; // @[StoreQueue.scala 250:20:@4837.4]
  assign io_storeAddrDone_14 = addrKnown_14; // @[StoreQueue.scala 250:20:@4838.4]
  assign io_storeAddrDone_15 = addrKnown_15; // @[StoreQueue.scala 250:20:@4839.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[StoreQueue.scala 249:20:@4808.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[StoreQueue.scala 249:20:@4809.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[StoreQueue.scala 249:20:@4810.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[StoreQueue.scala 249:20:@4811.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[StoreQueue.scala 249:20:@4812.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[StoreQueue.scala 249:20:@4813.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[StoreQueue.scala 249:20:@4814.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[StoreQueue.scala 249:20:@4815.4]
  assign io_storeDataDone_8 = dataKnown_8; // @[StoreQueue.scala 249:20:@4816.4]
  assign io_storeDataDone_9 = dataKnown_9; // @[StoreQueue.scala 249:20:@4817.4]
  assign io_storeDataDone_10 = dataKnown_10; // @[StoreQueue.scala 249:20:@4818.4]
  assign io_storeDataDone_11 = dataKnown_11; // @[StoreQueue.scala 249:20:@4819.4]
  assign io_storeDataDone_12 = dataKnown_12; // @[StoreQueue.scala 249:20:@4820.4]
  assign io_storeDataDone_13 = dataKnown_13; // @[StoreQueue.scala 249:20:@4821.4]
  assign io_storeDataDone_14 = dataKnown_14; // @[StoreQueue.scala 249:20:@4822.4]
  assign io_storeDataDone_15 = dataKnown_15; // @[StoreQueue.scala 249:20:@4823.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[StoreQueue.scala 247:21:@4776.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[StoreQueue.scala 247:21:@4777.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[StoreQueue.scala 247:21:@4778.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[StoreQueue.scala 247:21:@4779.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[StoreQueue.scala 247:21:@4780.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[StoreQueue.scala 247:21:@4781.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[StoreQueue.scala 247:21:@4782.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[StoreQueue.scala 247:21:@4783.4]
  assign io_storeAddrQueue_8 = addrQ_8; // @[StoreQueue.scala 247:21:@4784.4]
  assign io_storeAddrQueue_9 = addrQ_9; // @[StoreQueue.scala 247:21:@4785.4]
  assign io_storeAddrQueue_10 = addrQ_10; // @[StoreQueue.scala 247:21:@4786.4]
  assign io_storeAddrQueue_11 = addrQ_11; // @[StoreQueue.scala 247:21:@4787.4]
  assign io_storeAddrQueue_12 = addrQ_12; // @[StoreQueue.scala 247:21:@4788.4]
  assign io_storeAddrQueue_13 = addrQ_13; // @[StoreQueue.scala 247:21:@4789.4]
  assign io_storeAddrQueue_14 = addrQ_14; // @[StoreQueue.scala 247:21:@4790.4]
  assign io_storeAddrQueue_15 = addrQ_15; // @[StoreQueue.scala 247:21:@4791.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[StoreQueue.scala 248:21:@4792.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[StoreQueue.scala 248:21:@4793.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[StoreQueue.scala 248:21:@4794.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[StoreQueue.scala 248:21:@4795.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[StoreQueue.scala 248:21:@4796.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[StoreQueue.scala 248:21:@4797.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[StoreQueue.scala 248:21:@4798.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[StoreQueue.scala 248:21:@4799.4]
  assign io_storeDataQueue_8 = dataQ_8; // @[StoreQueue.scala 248:21:@4800.4]
  assign io_storeDataQueue_9 = dataQ_9; // @[StoreQueue.scala 248:21:@4801.4]
  assign io_storeDataQueue_10 = dataQ_10; // @[StoreQueue.scala 248:21:@4802.4]
  assign io_storeDataQueue_11 = dataQ_11; // @[StoreQueue.scala 248:21:@4803.4]
  assign io_storeDataQueue_12 = dataQ_12; // @[StoreQueue.scala 248:21:@4804.4]
  assign io_storeDataQueue_13 = dataQ_13; // @[StoreQueue.scala 248:21:@4805.4]
  assign io_storeDataQueue_14 = dataQ_14; // @[StoreQueue.scala 248:21:@4806.4]
  assign io_storeDataQueue_15 = dataQ_15; // @[StoreQueue.scala 248:21:@4807.4]
  assign io_storeAddrToMem = 4'hf == head ? addrQ_15 : _GEN_910; // @[StoreQueue.scala 253:21:@4842.4]
  assign io_storeDataToMem = 4'hf == head ? dataQ_15 : _GEN_1136; // @[StoreQueue.scala 252:21:@4841.4]
  assign io_storeEnableToMem = _T_3525 & _T_3542; // @[StoreQueue.scala 251:23:@4840.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  storeCompleted_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  storeCompleted_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  storeCompleted_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  storeCompleted_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  storeCompleted_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  storeCompleted_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  storeCompleted_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  storeCompleted_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  checkBits_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  checkBits_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  checkBits_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  checkBits_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  checkBits_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  checkBits_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  checkBits_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  checkBits_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  checkBits_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  checkBits_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  checkBits_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  checkBits_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  checkBits_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  checkBits_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  checkBits_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  checkBits_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  previousLoadHead = _RAND_146[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_1120[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_1121[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1804) begin
          offsetQ_0 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1804) begin
            offsetQ_0 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1804) begin
              offsetQ_0 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1804) begin
                offsetQ_0 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1804) begin
                  offsetQ_0 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1804) begin
                    offsetQ_0 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1804) begin
                      offsetQ_0 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1804) begin
                        offsetQ_0 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1804) begin
                          offsetQ_0 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1804) begin
                            offsetQ_0 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1804) begin
                              offsetQ_0 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1804) begin
                                offsetQ_0 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1804) begin
                                  offsetQ_0 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1804) begin
                                    offsetQ_0 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1804) begin
                                      offsetQ_0 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1822) begin
          offsetQ_1 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1822) begin
            offsetQ_1 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1822) begin
              offsetQ_1 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1822) begin
                offsetQ_1 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1822) begin
                  offsetQ_1 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1822) begin
                    offsetQ_1 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1822) begin
                      offsetQ_1 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1822) begin
                        offsetQ_1 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1822) begin
                          offsetQ_1 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1822) begin
                            offsetQ_1 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1822) begin
                              offsetQ_1 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1822) begin
                                offsetQ_1 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1822) begin
                                  offsetQ_1 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1822) begin
                                    offsetQ_1 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1822) begin
                                      offsetQ_1 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1840) begin
          offsetQ_2 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1840) begin
            offsetQ_2 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1840) begin
              offsetQ_2 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1840) begin
                offsetQ_2 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1840) begin
                  offsetQ_2 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1840) begin
                    offsetQ_2 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1840) begin
                      offsetQ_2 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1840) begin
                        offsetQ_2 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1840) begin
                          offsetQ_2 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1840) begin
                            offsetQ_2 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1840) begin
                              offsetQ_2 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1840) begin
                                offsetQ_2 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1840) begin
                                  offsetQ_2 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1840) begin
                                    offsetQ_2 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1840) begin
                                      offsetQ_2 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1858) begin
          offsetQ_3 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1858) begin
            offsetQ_3 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1858) begin
              offsetQ_3 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1858) begin
                offsetQ_3 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1858) begin
                  offsetQ_3 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1858) begin
                    offsetQ_3 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1858) begin
                      offsetQ_3 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1858) begin
                        offsetQ_3 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1858) begin
                          offsetQ_3 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1858) begin
                            offsetQ_3 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1858) begin
                              offsetQ_3 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1858) begin
                                offsetQ_3 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1858) begin
                                  offsetQ_3 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1858) begin
                                    offsetQ_3 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1858) begin
                                      offsetQ_3 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1876) begin
          offsetQ_4 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1876) begin
            offsetQ_4 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1876) begin
              offsetQ_4 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1876) begin
                offsetQ_4 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1876) begin
                  offsetQ_4 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1876) begin
                    offsetQ_4 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1876) begin
                      offsetQ_4 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1876) begin
                        offsetQ_4 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1876) begin
                          offsetQ_4 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1876) begin
                            offsetQ_4 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1876) begin
                              offsetQ_4 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1876) begin
                                offsetQ_4 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1876) begin
                                  offsetQ_4 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1876) begin
                                    offsetQ_4 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1876) begin
                                      offsetQ_4 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_1894) begin
          offsetQ_5 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1894) begin
            offsetQ_5 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1894) begin
              offsetQ_5 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1894) begin
                offsetQ_5 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1894) begin
                  offsetQ_5 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1894) begin
                    offsetQ_5 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1894) begin
                      offsetQ_5 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1894) begin
                        offsetQ_5 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1894) begin
                          offsetQ_5 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1894) begin
                            offsetQ_5 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1894) begin
                              offsetQ_5 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1894) begin
                                offsetQ_5 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1894) begin
                                  offsetQ_5 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1894) begin
                                    offsetQ_5 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1894) begin
                                      offsetQ_5 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_1912) begin
          offsetQ_6 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1912) begin
            offsetQ_6 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1912) begin
              offsetQ_6 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1912) begin
                offsetQ_6 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1912) begin
                  offsetQ_6 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1912) begin
                    offsetQ_6 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1912) begin
                      offsetQ_6 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1912) begin
                        offsetQ_6 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1912) begin
                          offsetQ_6 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1912) begin
                            offsetQ_6 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1912) begin
                              offsetQ_6 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1912) begin
                                offsetQ_6 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1912) begin
                                  offsetQ_6 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1912) begin
                                    offsetQ_6 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1912) begin
                                      offsetQ_6 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_1930) begin
          offsetQ_7 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1930) begin
            offsetQ_7 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1930) begin
              offsetQ_7 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1930) begin
                offsetQ_7 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1930) begin
                  offsetQ_7 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1930) begin
                    offsetQ_7 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1930) begin
                      offsetQ_7 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1930) begin
                        offsetQ_7 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1930) begin
                          offsetQ_7 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1930) begin
                            offsetQ_7 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1930) begin
                              offsetQ_7 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1930) begin
                                offsetQ_7 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1930) begin
                                  offsetQ_7 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1930) begin
                                    offsetQ_7 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1930) begin
                                      offsetQ_7 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_1948) begin
          offsetQ_8 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1948) begin
            offsetQ_8 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1948) begin
              offsetQ_8 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1948) begin
                offsetQ_8 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1948) begin
                  offsetQ_8 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1948) begin
                    offsetQ_8 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1948) begin
                      offsetQ_8 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1948) begin
                        offsetQ_8 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1948) begin
                          offsetQ_8 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1948) begin
                            offsetQ_8 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1948) begin
                              offsetQ_8 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1948) begin
                                offsetQ_8 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1948) begin
                                  offsetQ_8 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1948) begin
                                    offsetQ_8 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1948) begin
                                      offsetQ_8 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_1966) begin
          offsetQ_9 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1966) begin
            offsetQ_9 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1966) begin
              offsetQ_9 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1966) begin
                offsetQ_9 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1966) begin
                  offsetQ_9 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1966) begin
                    offsetQ_9 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1966) begin
                      offsetQ_9 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1966) begin
                        offsetQ_9 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1966) begin
                          offsetQ_9 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1966) begin
                            offsetQ_9 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1966) begin
                              offsetQ_9 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1966) begin
                                offsetQ_9 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1966) begin
                                  offsetQ_9 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1966) begin
                                    offsetQ_9 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1966) begin
                                      offsetQ_9 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_1984) begin
          offsetQ_10 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1984) begin
            offsetQ_10 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1984) begin
              offsetQ_10 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1984) begin
                offsetQ_10 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1984) begin
                  offsetQ_10 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1984) begin
                    offsetQ_10 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1984) begin
                      offsetQ_10 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1984) begin
                        offsetQ_10 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1984) begin
                          offsetQ_10 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1984) begin
                            offsetQ_10 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1984) begin
                              offsetQ_10 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1984) begin
                                offsetQ_10 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1984) begin
                                  offsetQ_10 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1984) begin
                                    offsetQ_10 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1984) begin
                                      offsetQ_10 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2002) begin
          offsetQ_11 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2002) begin
            offsetQ_11 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2002) begin
              offsetQ_11 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2002) begin
                offsetQ_11 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2002) begin
                  offsetQ_11 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2002) begin
                    offsetQ_11 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2002) begin
                      offsetQ_11 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2002) begin
                        offsetQ_11 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2002) begin
                          offsetQ_11 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2002) begin
                            offsetQ_11 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2002) begin
                              offsetQ_11 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2002) begin
                                offsetQ_11 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2002) begin
                                  offsetQ_11 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2002) begin
                                    offsetQ_11 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2002) begin
                                      offsetQ_11 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2020) begin
          offsetQ_12 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2020) begin
            offsetQ_12 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2020) begin
              offsetQ_12 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2020) begin
                offsetQ_12 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2020) begin
                  offsetQ_12 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2020) begin
                    offsetQ_12 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2020) begin
                      offsetQ_12 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2020) begin
                        offsetQ_12 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2020) begin
                          offsetQ_12 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2020) begin
                            offsetQ_12 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2020) begin
                              offsetQ_12 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2020) begin
                                offsetQ_12 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2020) begin
                                  offsetQ_12 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2020) begin
                                    offsetQ_12 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2020) begin
                                      offsetQ_12 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2038) begin
          offsetQ_13 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2038) begin
            offsetQ_13 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2038) begin
              offsetQ_13 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2038) begin
                offsetQ_13 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2038) begin
                  offsetQ_13 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2038) begin
                    offsetQ_13 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2038) begin
                      offsetQ_13 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2038) begin
                        offsetQ_13 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2038) begin
                          offsetQ_13 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2038) begin
                            offsetQ_13 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2038) begin
                              offsetQ_13 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2038) begin
                                offsetQ_13 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2038) begin
                                  offsetQ_13 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2038) begin
                                    offsetQ_13 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2038) begin
                                      offsetQ_13 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2056) begin
          offsetQ_14 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2056) begin
            offsetQ_14 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2056) begin
              offsetQ_14 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2056) begin
                offsetQ_14 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2056) begin
                  offsetQ_14 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2056) begin
                    offsetQ_14 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2056) begin
                      offsetQ_14 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2056) begin
                        offsetQ_14 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2056) begin
                          offsetQ_14 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2056) begin
                            offsetQ_14 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2056) begin
                              offsetQ_14 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2056) begin
                                offsetQ_14 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2056) begin
                                  offsetQ_14 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2056) begin
                                    offsetQ_14 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2056) begin
                                      offsetQ_14 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2074) begin
          offsetQ_15 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2074) begin
            offsetQ_15 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2074) begin
              offsetQ_15 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2074) begin
                offsetQ_15 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2074) begin
                  offsetQ_15 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2074) begin
                    offsetQ_15 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2074) begin
                      offsetQ_15 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2074) begin
                        offsetQ_15 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2074) begin
                          offsetQ_15 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2074) begin
                            offsetQ_15 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2074) begin
                              offsetQ_15 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2074) begin
                                offsetQ_15 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2074) begin
                                  offsetQ_15 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2074) begin
                                    offsetQ_15 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2074) begin
                                      offsetQ_15 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7582) begin
          addrQ_0 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7618) begin
          addrQ_1 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7654) begin
          addrQ_2 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7690) begin
          addrQ_3 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7726) begin
          addrQ_4 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7762) begin
          addrQ_5 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7798) begin
          addrQ_6 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7834) begin
          addrQ_7 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7870) begin
          addrQ_8 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7906) begin
          addrQ_9 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7942) begin
          addrQ_10 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7978) begin
          addrQ_11 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8014) begin
          addrQ_12 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8050) begin
          addrQ_13 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8086) begin
          addrQ_14 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8122) begin
          addrQ_15 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7599) begin
          dataQ_0 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7635) begin
          dataQ_1 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7671) begin
          dataQ_2 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7707) begin
          dataQ_3 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7743) begin
          dataQ_4 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7779) begin
          dataQ_5 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7815) begin
          dataQ_6 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7851) begin
          dataQ_7 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7887) begin
          dataQ_8 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7923) begin
          dataQ_9 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7959) begin
          dataQ_10 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7995) begin
          dataQ_11 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8031) begin
          dataQ_12 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8067) begin
          dataQ_13 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8103) begin
          dataQ_14 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8139) begin
          dataQ_15 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_7582) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_7618) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_7654) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_7690) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_7726) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_7762) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_7798) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_7834) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_7870) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_7906) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_7942) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_7978) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_8014) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_8050) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_8086) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_8122) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_7599) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_7635) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_7671) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_7707) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_7743) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_7779) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_7815) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_7851) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_7887) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_7923) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_7959) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_7995) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_8031) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_8067) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_8103) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_8139) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1758;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1759;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1760;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1761;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1762;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1763;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1764;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1765;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1766;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1767;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1768;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1769;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1770;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1771;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1772;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1773;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_3547) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_3553) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_3559) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_3565) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_3571) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_3577) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_3583) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_3589) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        storeCompleted_8 <= 1'h0;
      end else begin
        if (_T_3595) begin
          storeCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        storeCompleted_9 <= 1'h0;
      end else begin
        if (_T_3601) begin
          storeCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        storeCompleted_10 <= 1'h0;
      end else begin
        if (_T_3607) begin
          storeCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        storeCompleted_11 <= 1'h0;
      end else begin
        if (_T_3613) begin
          storeCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        storeCompleted_12 <= 1'h0;
      end else begin
        if (_T_3619) begin
          storeCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        storeCompleted_13 <= 1'h0;
      end else begin
        if (_T_3625) begin
          storeCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        storeCompleted_14 <= 1'h0;
      end else begin
        if (_T_3631) begin
          storeCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        storeCompleted_15 <= 1'h0;
      end else begin
        if (_T_3637) begin
          storeCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2101;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2105) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2113) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2131;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2135) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2143) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2161;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2165) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2173) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2191;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2195) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2203) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2221;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2225) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2233) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2251;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2255) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2263) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2281;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2285) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2293) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2311;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2315) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2323) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2341;
      end else begin
        if (io_loadEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2345) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2353) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2371;
      end else begin
        if (io_loadEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2375) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2383) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2401;
      end else begin
        if (io_loadEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2405) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2413) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2431;
      end else begin
        if (io_loadEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2435) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2443) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2461;
      end else begin
        if (io_loadEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2465) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2473) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2491;
      end else begin
        if (io_loadEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2495) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2503) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2521;
      end else begin
        if (io_loadEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2525) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2533) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2551;
      end else begin
        if (io_loadEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2555) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2563) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_A( // @[:@4844.2]
  input         clock, // @[:@4845.4]
  input         reset, // @[:@4846.4]
  input         io_bbStart, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_0, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_1, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_2, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_3, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_4, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_5, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_6, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_7, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_8, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_9, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_10, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_11, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_12, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_13, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_14, // @[:@4847.4]
  input  [3:0]  io_bbLoadOffsets_15, // @[:@4847.4]
  input         io_bbNumLoads, // @[:@4847.4]
  output [3:0]  io_loadTail, // @[:@4847.4]
  output [3:0]  io_loadHead, // @[:@4847.4]
  output        io_loadEmpty, // @[:@4847.4]
  input  [3:0]  io_storeTail, // @[:@4847.4]
  input  [3:0]  io_storeHead, // @[:@4847.4]
  input         io_storeEmpty, // @[:@4847.4]
  input         io_storeAddrDone_0, // @[:@4847.4]
  input         io_storeAddrDone_1, // @[:@4847.4]
  input         io_storeAddrDone_2, // @[:@4847.4]
  input         io_storeAddrDone_3, // @[:@4847.4]
  input         io_storeAddrDone_4, // @[:@4847.4]
  input         io_storeAddrDone_5, // @[:@4847.4]
  input         io_storeAddrDone_6, // @[:@4847.4]
  input         io_storeAddrDone_7, // @[:@4847.4]
  input         io_storeAddrDone_8, // @[:@4847.4]
  input         io_storeAddrDone_9, // @[:@4847.4]
  input         io_storeAddrDone_10, // @[:@4847.4]
  input         io_storeAddrDone_11, // @[:@4847.4]
  input         io_storeAddrDone_12, // @[:@4847.4]
  input         io_storeAddrDone_13, // @[:@4847.4]
  input         io_storeAddrDone_14, // @[:@4847.4]
  input         io_storeAddrDone_15, // @[:@4847.4]
  input         io_storeDataDone_0, // @[:@4847.4]
  input         io_storeDataDone_1, // @[:@4847.4]
  input         io_storeDataDone_2, // @[:@4847.4]
  input         io_storeDataDone_3, // @[:@4847.4]
  input         io_storeDataDone_4, // @[:@4847.4]
  input         io_storeDataDone_5, // @[:@4847.4]
  input         io_storeDataDone_6, // @[:@4847.4]
  input         io_storeDataDone_7, // @[:@4847.4]
  input         io_storeDataDone_8, // @[:@4847.4]
  input         io_storeDataDone_9, // @[:@4847.4]
  input         io_storeDataDone_10, // @[:@4847.4]
  input         io_storeDataDone_11, // @[:@4847.4]
  input         io_storeDataDone_12, // @[:@4847.4]
  input         io_storeDataDone_13, // @[:@4847.4]
  input         io_storeDataDone_14, // @[:@4847.4]
  input         io_storeDataDone_15, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_0, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_1, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_2, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_3, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_4, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_5, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_6, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_7, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_8, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_9, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_10, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_11, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_12, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_13, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_14, // @[:@4847.4]
  input  [31:0] io_storeAddrQueue_15, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_0, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_1, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_2, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_3, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_4, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_5, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_6, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_7, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_8, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_9, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_10, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_11, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_12, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_13, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_14, // @[:@4847.4]
  input  [31:0] io_storeDataQueue_15, // @[:@4847.4]
  output        io_loadAddrDone_0, // @[:@4847.4]
  output        io_loadAddrDone_1, // @[:@4847.4]
  output        io_loadAddrDone_2, // @[:@4847.4]
  output        io_loadAddrDone_3, // @[:@4847.4]
  output        io_loadAddrDone_4, // @[:@4847.4]
  output        io_loadAddrDone_5, // @[:@4847.4]
  output        io_loadAddrDone_6, // @[:@4847.4]
  output        io_loadAddrDone_7, // @[:@4847.4]
  output        io_loadAddrDone_8, // @[:@4847.4]
  output        io_loadAddrDone_9, // @[:@4847.4]
  output        io_loadAddrDone_10, // @[:@4847.4]
  output        io_loadAddrDone_11, // @[:@4847.4]
  output        io_loadAddrDone_12, // @[:@4847.4]
  output        io_loadAddrDone_13, // @[:@4847.4]
  output        io_loadAddrDone_14, // @[:@4847.4]
  output        io_loadAddrDone_15, // @[:@4847.4]
  output        io_loadDataDone_0, // @[:@4847.4]
  output        io_loadDataDone_1, // @[:@4847.4]
  output        io_loadDataDone_2, // @[:@4847.4]
  output        io_loadDataDone_3, // @[:@4847.4]
  output        io_loadDataDone_4, // @[:@4847.4]
  output        io_loadDataDone_5, // @[:@4847.4]
  output        io_loadDataDone_6, // @[:@4847.4]
  output        io_loadDataDone_7, // @[:@4847.4]
  output        io_loadDataDone_8, // @[:@4847.4]
  output        io_loadDataDone_9, // @[:@4847.4]
  output        io_loadDataDone_10, // @[:@4847.4]
  output        io_loadDataDone_11, // @[:@4847.4]
  output        io_loadDataDone_12, // @[:@4847.4]
  output        io_loadDataDone_13, // @[:@4847.4]
  output        io_loadDataDone_14, // @[:@4847.4]
  output        io_loadDataDone_15, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_0, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_1, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_2, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_3, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_4, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_5, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_6, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_7, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_8, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_9, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_10, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_11, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_12, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_13, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_14, // @[:@4847.4]
  output [31:0] io_loadAddrQueue_15, // @[:@4847.4]
  input         io_loadAddrEnable_0, // @[:@4847.4]
  input  [31:0] io_addrFromLoadPorts_0, // @[:@4847.4]
  input         io_loadPorts_0_ready, // @[:@4847.4]
  output        io_loadPorts_0_valid, // @[:@4847.4]
  output [31:0] io_loadPorts_0_bits, // @[:@4847.4]
  input  [31:0] io_loadDataFromMem, // @[:@4847.4]
  output [31:0] io_loadAddrToMem, // @[:@4847.4]
  output        io_loadEnableToMem, // @[:@4847.4]
  input         io_memIsReadyForLoads // @[:@4847.4]
);
  reg [3:0] head; // @[LoadQueue.scala 50:21:@4849.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[LoadQueue.scala 51:21:@4850.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[LoadQueue.scala 53:24:@4868.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[LoadQueue.scala 54:22:@4886.4]
  reg [31:0] _RAND_33;
  reg [31:0] addrQ_0; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_34;
  reg [31:0] addrQ_1; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_35;
  reg [31:0] addrQ_2; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_36;
  reg [31:0] addrQ_3; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_37;
  reg [31:0] addrQ_4; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_38;
  reg [31:0] addrQ_5; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_39;
  reg [31:0] addrQ_6; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_40;
  reg [31:0] addrQ_7; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_41;
  reg [31:0] addrQ_8; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_42;
  reg [31:0] addrQ_9; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_43;
  reg [31:0] addrQ_10; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_44;
  reg [31:0] addrQ_11; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_45;
  reg [31:0] addrQ_12; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_46;
  reg [31:0] addrQ_13; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_47;
  reg [31:0] addrQ_14; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_48;
  reg [31:0] addrQ_15; // @[LoadQueue.scala 55:22:@4904.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[LoadQueue.scala 56:22:@4922.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[LoadQueue.scala 57:26:@4940.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[LoadQueue.scala 58:26:@4958.4]
  reg [31:0] _RAND_97;
  reg  loadCompleted_0; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_98;
  reg  loadCompleted_1; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_99;
  reg  loadCompleted_2; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_100;
  reg  loadCompleted_3; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_101;
  reg  loadCompleted_4; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_102;
  reg  loadCompleted_5; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_103;
  reg  loadCompleted_6; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_104;
  reg  loadCompleted_7; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_105;
  reg  loadCompleted_8; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_106;
  reg  loadCompleted_9; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_107;
  reg  loadCompleted_10; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_108;
  reg  loadCompleted_11; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_109;
  reg  loadCompleted_12; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_110;
  reg  loadCompleted_13; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_111;
  reg  loadCompleted_14; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_112;
  reg  loadCompleted_15; // @[LoadQueue.scala 59:30:@4976.4]
  reg [31:0] _RAND_113;
  reg  allocatedEntries_0; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_114;
  reg  allocatedEntries_1; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_115;
  reg  allocatedEntries_2; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_116;
  reg  allocatedEntries_3; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_117;
  reg  allocatedEntries_4; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_118;
  reg  allocatedEntries_5; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_119;
  reg  allocatedEntries_6; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_120;
  reg  allocatedEntries_7; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_121;
  reg  allocatedEntries_8; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_122;
  reg  allocatedEntries_9; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_123;
  reg  allocatedEntries_10; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_124;
  reg  allocatedEntries_11; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_125;
  reg  allocatedEntries_12; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_126;
  reg  allocatedEntries_13; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_127;
  reg  allocatedEntries_14; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_128;
  reg  allocatedEntries_15; // @[LoadQueue.scala 60:33:@4994.4]
  reg [31:0] _RAND_129;
  reg  bypassInitiated_0; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_130;
  reg  bypassInitiated_1; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_131;
  reg  bypassInitiated_2; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_132;
  reg  bypassInitiated_3; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_133;
  reg  bypassInitiated_4; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_134;
  reg  bypassInitiated_5; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_135;
  reg  bypassInitiated_6; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_136;
  reg  bypassInitiated_7; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_137;
  reg  bypassInitiated_8; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_138;
  reg  bypassInitiated_9; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_139;
  reg  bypassInitiated_10; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_140;
  reg  bypassInitiated_11; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_141;
  reg  bypassInitiated_12; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_142;
  reg  bypassInitiated_13; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_143;
  reg  bypassInitiated_14; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_144;
  reg  bypassInitiated_15; // @[LoadQueue.scala 61:32:@5012.4]
  reg [31:0] _RAND_145;
  reg  checkBits_0; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_146;
  reg  checkBits_1; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_147;
  reg  checkBits_2; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_148;
  reg  checkBits_3; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_149;
  reg  checkBits_4; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_150;
  reg  checkBits_5; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_151;
  reg  checkBits_6; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_152;
  reg  checkBits_7; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_153;
  reg  checkBits_8; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_154;
  reg  checkBits_9; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_155;
  reg  checkBits_10; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_156;
  reg  checkBits_11; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_157;
  reg  checkBits_12; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_158;
  reg  checkBits_13; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_159;
  reg  checkBits_14; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_160;
  reg  checkBits_15; // @[LoadQueue.scala 62:26:@5030.4]
  reg [31:0] _RAND_161;
  wire [5:0] _GEN_2262; // @[util.scala 14:20:@5032.4]
  wire [6:0] _T_1716; // @[util.scala 14:20:@5032.4]
  wire [6:0] _T_1717; // @[util.scala 14:20:@5033.4]
  wire [5:0] _T_1718; // @[util.scala 14:20:@5034.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@5035.4]
  wire [4:0] _T_1719; // @[util.scala 14:25:@5035.4]
  wire [4:0] _GEN_2263; // @[LoadQueue.scala 71:46:@5036.4]
  wire  _T_1720; // @[LoadQueue.scala 71:46:@5036.4]
  wire  initBits_0; // @[LoadQueue.scala 71:63:@5037.4]
  wire [6:0] _T_1725; // @[util.scala 14:20:@5039.4]
  wire [6:0] _T_1726; // @[util.scala 14:20:@5040.4]
  wire [5:0] _T_1727; // @[util.scala 14:20:@5041.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@5042.4]
  wire [4:0] _T_1728; // @[util.scala 14:25:@5042.4]
  wire  _T_1729; // @[LoadQueue.scala 71:46:@5043.4]
  wire  initBits_1; // @[LoadQueue.scala 71:63:@5044.4]
  wire [6:0] _T_1734; // @[util.scala 14:20:@5046.4]
  wire [6:0] _T_1735; // @[util.scala 14:20:@5047.4]
  wire [5:0] _T_1736; // @[util.scala 14:20:@5048.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@5049.4]
  wire [4:0] _T_1737; // @[util.scala 14:25:@5049.4]
  wire  _T_1738; // @[LoadQueue.scala 71:46:@5050.4]
  wire  initBits_2; // @[LoadQueue.scala 71:63:@5051.4]
  wire [6:0] _T_1743; // @[util.scala 14:20:@5053.4]
  wire [6:0] _T_1744; // @[util.scala 14:20:@5054.4]
  wire [5:0] _T_1745; // @[util.scala 14:20:@5055.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@5056.4]
  wire [4:0] _T_1746; // @[util.scala 14:25:@5056.4]
  wire  _T_1747; // @[LoadQueue.scala 71:46:@5057.4]
  wire  initBits_3; // @[LoadQueue.scala 71:63:@5058.4]
  wire [6:0] _T_1752; // @[util.scala 14:20:@5060.4]
  wire [6:0] _T_1753; // @[util.scala 14:20:@5061.4]
  wire [5:0] _T_1754; // @[util.scala 14:20:@5062.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@5063.4]
  wire [4:0] _T_1755; // @[util.scala 14:25:@5063.4]
  wire  _T_1756; // @[LoadQueue.scala 71:46:@5064.4]
  wire  initBits_4; // @[LoadQueue.scala 71:63:@5065.4]
  wire [6:0] _T_1761; // @[util.scala 14:20:@5067.4]
  wire [6:0] _T_1762; // @[util.scala 14:20:@5068.4]
  wire [5:0] _T_1763; // @[util.scala 14:20:@5069.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@5070.4]
  wire [4:0] _T_1764; // @[util.scala 14:25:@5070.4]
  wire  _T_1765; // @[LoadQueue.scala 71:46:@5071.4]
  wire  initBits_5; // @[LoadQueue.scala 71:63:@5072.4]
  wire [6:0] _T_1770; // @[util.scala 14:20:@5074.4]
  wire [6:0] _T_1771; // @[util.scala 14:20:@5075.4]
  wire [5:0] _T_1772; // @[util.scala 14:20:@5076.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@5077.4]
  wire [4:0] _T_1773; // @[util.scala 14:25:@5077.4]
  wire  _T_1774; // @[LoadQueue.scala 71:46:@5078.4]
  wire  initBits_6; // @[LoadQueue.scala 71:63:@5079.4]
  wire [6:0] _T_1779; // @[util.scala 14:20:@5081.4]
  wire [6:0] _T_1780; // @[util.scala 14:20:@5082.4]
  wire [5:0] _T_1781; // @[util.scala 14:20:@5083.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@5084.4]
  wire [4:0] _T_1782; // @[util.scala 14:25:@5084.4]
  wire  _T_1783; // @[LoadQueue.scala 71:46:@5085.4]
  wire  initBits_7; // @[LoadQueue.scala 71:63:@5086.4]
  wire [6:0] _T_1788; // @[util.scala 14:20:@5088.4]
  wire [6:0] _T_1789; // @[util.scala 14:20:@5089.4]
  wire [5:0] _T_1790; // @[util.scala 14:20:@5090.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@5091.4]
  wire [4:0] _T_1791; // @[util.scala 14:25:@5091.4]
  wire  _T_1792; // @[LoadQueue.scala 71:46:@5092.4]
  wire  initBits_8; // @[LoadQueue.scala 71:63:@5093.4]
  wire [6:0] _T_1797; // @[util.scala 14:20:@5095.4]
  wire [6:0] _T_1798; // @[util.scala 14:20:@5096.4]
  wire [5:0] _T_1799; // @[util.scala 14:20:@5097.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@5098.4]
  wire [4:0] _T_1800; // @[util.scala 14:25:@5098.4]
  wire  _T_1801; // @[LoadQueue.scala 71:46:@5099.4]
  wire  initBits_9; // @[LoadQueue.scala 71:63:@5100.4]
  wire [6:0] _T_1806; // @[util.scala 14:20:@5102.4]
  wire [6:0] _T_1807; // @[util.scala 14:20:@5103.4]
  wire [5:0] _T_1808; // @[util.scala 14:20:@5104.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@5105.4]
  wire [4:0] _T_1809; // @[util.scala 14:25:@5105.4]
  wire  _T_1810; // @[LoadQueue.scala 71:46:@5106.4]
  wire  initBits_10; // @[LoadQueue.scala 71:63:@5107.4]
  wire [6:0] _T_1815; // @[util.scala 14:20:@5109.4]
  wire [6:0] _T_1816; // @[util.scala 14:20:@5110.4]
  wire [5:0] _T_1817; // @[util.scala 14:20:@5111.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@5112.4]
  wire [4:0] _T_1818; // @[util.scala 14:25:@5112.4]
  wire  _T_1819; // @[LoadQueue.scala 71:46:@5113.4]
  wire  initBits_11; // @[LoadQueue.scala 71:63:@5114.4]
  wire [6:0] _T_1824; // @[util.scala 14:20:@5116.4]
  wire [6:0] _T_1825; // @[util.scala 14:20:@5117.4]
  wire [5:0] _T_1826; // @[util.scala 14:20:@5118.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@5119.4]
  wire [4:0] _T_1827; // @[util.scala 14:25:@5119.4]
  wire  _T_1828; // @[LoadQueue.scala 71:46:@5120.4]
  wire  initBits_12; // @[LoadQueue.scala 71:63:@5121.4]
  wire [6:0] _T_1833; // @[util.scala 14:20:@5123.4]
  wire [6:0] _T_1834; // @[util.scala 14:20:@5124.4]
  wire [5:0] _T_1835; // @[util.scala 14:20:@5125.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@5126.4]
  wire [4:0] _T_1836; // @[util.scala 14:25:@5126.4]
  wire  _T_1837; // @[LoadQueue.scala 71:46:@5127.4]
  wire  initBits_13; // @[LoadQueue.scala 71:63:@5128.4]
  wire [6:0] _T_1842; // @[util.scala 14:20:@5130.4]
  wire [6:0] _T_1843; // @[util.scala 14:20:@5131.4]
  wire [5:0] _T_1844; // @[util.scala 14:20:@5132.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@5133.4]
  wire [4:0] _T_1845; // @[util.scala 14:25:@5133.4]
  wire  _T_1846; // @[LoadQueue.scala 71:46:@5134.4]
  wire  initBits_14; // @[LoadQueue.scala 71:63:@5135.4]
  wire [6:0] _T_1851; // @[util.scala 14:20:@5137.4]
  wire [6:0] _T_1852; // @[util.scala 14:20:@5138.4]
  wire [5:0] _T_1853; // @[util.scala 14:20:@5139.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@5140.4]
  wire [4:0] _T_1854; // @[util.scala 14:25:@5140.4]
  wire  _T_1855; // @[LoadQueue.scala 71:46:@5141.4]
  wire  initBits_15; // @[LoadQueue.scala 71:63:@5142.4]
  wire  _T_1878; // @[LoadQueue.scala 73:78:@5160.4]
  wire  _T_1879; // @[LoadQueue.scala 73:78:@5161.4]
  wire  _T_1880; // @[LoadQueue.scala 73:78:@5162.4]
  wire  _T_1881; // @[LoadQueue.scala 73:78:@5163.4]
  wire  _T_1882; // @[LoadQueue.scala 73:78:@5164.4]
  wire  _T_1883; // @[LoadQueue.scala 73:78:@5165.4]
  wire  _T_1884; // @[LoadQueue.scala 73:78:@5166.4]
  wire  _T_1885; // @[LoadQueue.scala 73:78:@5167.4]
  wire  _T_1886; // @[LoadQueue.scala 73:78:@5168.4]
  wire  _T_1887; // @[LoadQueue.scala 73:78:@5169.4]
  wire  _T_1888; // @[LoadQueue.scala 73:78:@5170.4]
  wire  _T_1889; // @[LoadQueue.scala 73:78:@5171.4]
  wire  _T_1890; // @[LoadQueue.scala 73:78:@5172.4]
  wire  _T_1891; // @[LoadQueue.scala 73:78:@5173.4]
  wire  _T_1892; // @[LoadQueue.scala 73:78:@5174.4]
  wire  _T_1893; // @[LoadQueue.scala 73:78:@5175.4]
  wire [3:0] _T_1924; // @[:@5215.6]
  wire [3:0] _GEN_1; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_2; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_3; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_4; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_5; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_6; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_7; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_8; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_9; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_10; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_11; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_12; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_13; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_14; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_15; // @[LoadQueue.scala 77:20:@5216.6]
  wire [3:0] _GEN_32; // @[LoadQueue.scala 76:25:@5209.4]
  wire  _GEN_33; // @[LoadQueue.scala 76:25:@5209.4]
  wire [3:0] _T_1942; // @[:@5231.6]
  wire [3:0] _GEN_35; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_36; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_37; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_38; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_39; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_40; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_41; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_42; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_43; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_44; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_45; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_46; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_47; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_48; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_49; // @[LoadQueue.scala 77:20:@5232.6]
  wire [3:0] _GEN_66; // @[LoadQueue.scala 76:25:@5225.4]
  wire  _GEN_67; // @[LoadQueue.scala 76:25:@5225.4]
  wire [3:0] _T_1960; // @[:@5247.6]
  wire [3:0] _GEN_69; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_70; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_71; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_72; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_73; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_74; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_75; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_76; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_77; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_78; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_79; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_80; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_81; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_82; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_83; // @[LoadQueue.scala 77:20:@5248.6]
  wire [3:0] _GEN_100; // @[LoadQueue.scala 76:25:@5241.4]
  wire  _GEN_101; // @[LoadQueue.scala 76:25:@5241.4]
  wire [3:0] _T_1978; // @[:@5263.6]
  wire [3:0] _GEN_103; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_104; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_105; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_106; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_107; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_108; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_109; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_110; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_111; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_112; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_113; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_114; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_115; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_116; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_117; // @[LoadQueue.scala 77:20:@5264.6]
  wire [3:0] _GEN_134; // @[LoadQueue.scala 76:25:@5257.4]
  wire  _GEN_135; // @[LoadQueue.scala 76:25:@5257.4]
  wire [3:0] _T_1996; // @[:@5279.6]
  wire [3:0] _GEN_137; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_138; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_139; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_140; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_141; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_142; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_143; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_144; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_145; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_146; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_147; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_148; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_149; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_150; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_151; // @[LoadQueue.scala 77:20:@5280.6]
  wire [3:0] _GEN_168; // @[LoadQueue.scala 76:25:@5273.4]
  wire  _GEN_169; // @[LoadQueue.scala 76:25:@5273.4]
  wire [3:0] _T_2014; // @[:@5295.6]
  wire [3:0] _GEN_171; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_172; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_173; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_174; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_175; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_176; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_177; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_178; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_179; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_180; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_181; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_182; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_183; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_184; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_185; // @[LoadQueue.scala 77:20:@5296.6]
  wire [3:0] _GEN_202; // @[LoadQueue.scala 76:25:@5289.4]
  wire  _GEN_203; // @[LoadQueue.scala 76:25:@5289.4]
  wire [3:0] _T_2032; // @[:@5311.6]
  wire [3:0] _GEN_205; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_206; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_207; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_208; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_209; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_210; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_211; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_212; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_213; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_214; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_215; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_216; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_217; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_218; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_219; // @[LoadQueue.scala 77:20:@5312.6]
  wire [3:0] _GEN_236; // @[LoadQueue.scala 76:25:@5305.4]
  wire  _GEN_237; // @[LoadQueue.scala 76:25:@5305.4]
  wire [3:0] _T_2050; // @[:@5327.6]
  wire [3:0] _GEN_239; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_240; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_241; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_242; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_243; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_244; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_245; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_246; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_247; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_248; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_249; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_250; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_251; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_252; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_253; // @[LoadQueue.scala 77:20:@5328.6]
  wire [3:0] _GEN_270; // @[LoadQueue.scala 76:25:@5321.4]
  wire  _GEN_271; // @[LoadQueue.scala 76:25:@5321.4]
  wire [3:0] _T_2068; // @[:@5343.6]
  wire [3:0] _GEN_273; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_274; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_275; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_276; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_277; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_278; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_279; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_280; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_281; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_282; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_283; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_284; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_285; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_286; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_287; // @[LoadQueue.scala 77:20:@5344.6]
  wire [3:0] _GEN_304; // @[LoadQueue.scala 76:25:@5337.4]
  wire  _GEN_305; // @[LoadQueue.scala 76:25:@5337.4]
  wire [3:0] _T_2086; // @[:@5359.6]
  wire [3:0] _GEN_307; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_308; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_309; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_310; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_311; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_312; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_313; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_314; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_315; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_316; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_317; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_318; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_319; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_320; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_321; // @[LoadQueue.scala 77:20:@5360.6]
  wire [3:0] _GEN_338; // @[LoadQueue.scala 76:25:@5353.4]
  wire  _GEN_339; // @[LoadQueue.scala 76:25:@5353.4]
  wire [3:0] _T_2104; // @[:@5375.6]
  wire [3:0] _GEN_341; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_342; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_343; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_344; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_345; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_346; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_347; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_348; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_349; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_350; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_351; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_352; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_353; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_354; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_355; // @[LoadQueue.scala 77:20:@5376.6]
  wire [3:0] _GEN_372; // @[LoadQueue.scala 76:25:@5369.4]
  wire  _GEN_373; // @[LoadQueue.scala 76:25:@5369.4]
  wire [3:0] _T_2122; // @[:@5391.6]
  wire [3:0] _GEN_375; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_376; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_377; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_378; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_379; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_380; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_381; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_382; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_383; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_384; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_385; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_386; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_387; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_388; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_389; // @[LoadQueue.scala 77:20:@5392.6]
  wire [3:0] _GEN_406; // @[LoadQueue.scala 76:25:@5385.4]
  wire  _GEN_407; // @[LoadQueue.scala 76:25:@5385.4]
  wire [3:0] _T_2140; // @[:@5407.6]
  wire [3:0] _GEN_409; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_410; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_411; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_412; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_413; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_414; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_415; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_416; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_417; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_418; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_419; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_420; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_421; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_422; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_423; // @[LoadQueue.scala 77:20:@5408.6]
  wire [3:0] _GEN_440; // @[LoadQueue.scala 76:25:@5401.4]
  wire  _GEN_441; // @[LoadQueue.scala 76:25:@5401.4]
  wire [3:0] _T_2158; // @[:@5423.6]
  wire [3:0] _GEN_443; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_444; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_445; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_446; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_447; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_448; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_449; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_450; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_451; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_452; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_453; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_454; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_455; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_456; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_457; // @[LoadQueue.scala 77:20:@5424.6]
  wire [3:0] _GEN_474; // @[LoadQueue.scala 76:25:@5417.4]
  wire  _GEN_475; // @[LoadQueue.scala 76:25:@5417.4]
  wire [3:0] _T_2176; // @[:@5439.6]
  wire [3:0] _GEN_477; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_478; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_479; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_480; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_481; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_482; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_483; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_484; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_485; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_486; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_487; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_488; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_489; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_490; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_491; // @[LoadQueue.scala 77:20:@5440.6]
  wire [3:0] _GEN_508; // @[LoadQueue.scala 76:25:@5433.4]
  wire  _GEN_509; // @[LoadQueue.scala 76:25:@5433.4]
  wire [3:0] _T_2194; // @[:@5455.6]
  wire [3:0] _GEN_511; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_512; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_513; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_514; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_515; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_516; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_517; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_518; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_519; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_520; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_521; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_522; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_523; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_524; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_525; // @[LoadQueue.scala 77:20:@5456.6]
  wire [3:0] _GEN_542; // @[LoadQueue.scala 76:25:@5449.4]
  wire  _GEN_543; // @[LoadQueue.scala 76:25:@5449.4]
  reg [3:0] previousStoreHead; // @[LoadQueue.scala 93:34:@5465.4]
  reg [31:0] _RAND_162;
  wire [4:0] _T_2216; // @[util.scala 10:8:@5474.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@5475.6]
  wire [4:0] _T_2217; // @[util.scala 10:14:@5475.6]
  wire [4:0] _GEN_2327; // @[LoadQueue.scala 97:56:@5476.6]
  wire  _T_2218; // @[LoadQueue.scala 97:56:@5476.6]
  wire  _T_2219; // @[LoadQueue.scala 96:50:@5477.6]
  wire  _T_2221; // @[LoadQueue.scala 96:34:@5478.6]
  wire  _T_2223; // @[LoadQueue.scala 101:36:@5486.8]
  wire  _T_2224; // @[LoadQueue.scala 101:86:@5487.8]
  wire  _T_2225; // @[LoadQueue.scala 101:61:@5488.8]
  wire  _T_2227; // @[LoadQueue.scala 103:36:@5493.10]
  wire  _T_2228; // @[LoadQueue.scala 103:69:@5494.10]
  wire  _T_2229; // @[LoadQueue.scala 104:31:@5495.10]
  wire  _T_2230; // @[LoadQueue.scala 103:94:@5496.10]
  wire  _T_2232; // @[LoadQueue.scala 103:54:@5497.10]
  wire  _T_2233; // @[LoadQueue.scala 103:51:@5498.10]
  wire  _GEN_560; // @[LoadQueue.scala 104:53:@5499.10]
  wire  _GEN_561; // @[LoadQueue.scala 101:102:@5489.8]
  wire  _GEN_562; // @[LoadQueue.scala 99:27:@5482.6]
  wire  _GEN_563; // @[LoadQueue.scala 95:34:@5467.4]
  wire [4:0] _T_2246; // @[util.scala 10:8:@5510.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@5511.6]
  wire [4:0] _T_2247; // @[util.scala 10:14:@5511.6]
  wire  _T_2248; // @[LoadQueue.scala 97:56:@5512.6]
  wire  _T_2249; // @[LoadQueue.scala 96:50:@5513.6]
  wire  _T_2251; // @[LoadQueue.scala 96:34:@5514.6]
  wire  _T_2253; // @[LoadQueue.scala 101:36:@5522.8]
  wire  _T_2254; // @[LoadQueue.scala 101:86:@5523.8]
  wire  _T_2255; // @[LoadQueue.scala 101:61:@5524.8]
  wire  _T_2258; // @[LoadQueue.scala 103:69:@5530.10]
  wire  _T_2259; // @[LoadQueue.scala 104:31:@5531.10]
  wire  _T_2260; // @[LoadQueue.scala 103:94:@5532.10]
  wire  _T_2262; // @[LoadQueue.scala 103:54:@5533.10]
  wire  _T_2263; // @[LoadQueue.scala 103:51:@5534.10]
  wire  _GEN_580; // @[LoadQueue.scala 104:53:@5535.10]
  wire  _GEN_581; // @[LoadQueue.scala 101:102:@5525.8]
  wire  _GEN_582; // @[LoadQueue.scala 99:27:@5518.6]
  wire  _GEN_583; // @[LoadQueue.scala 95:34:@5503.4]
  wire [4:0] _T_2276; // @[util.scala 10:8:@5546.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@5547.6]
  wire [4:0] _T_2277; // @[util.scala 10:14:@5547.6]
  wire  _T_2278; // @[LoadQueue.scala 97:56:@5548.6]
  wire  _T_2279; // @[LoadQueue.scala 96:50:@5549.6]
  wire  _T_2281; // @[LoadQueue.scala 96:34:@5550.6]
  wire  _T_2283; // @[LoadQueue.scala 101:36:@5558.8]
  wire  _T_2284; // @[LoadQueue.scala 101:86:@5559.8]
  wire  _T_2285; // @[LoadQueue.scala 101:61:@5560.8]
  wire  _T_2288; // @[LoadQueue.scala 103:69:@5566.10]
  wire  _T_2289; // @[LoadQueue.scala 104:31:@5567.10]
  wire  _T_2290; // @[LoadQueue.scala 103:94:@5568.10]
  wire  _T_2292; // @[LoadQueue.scala 103:54:@5569.10]
  wire  _T_2293; // @[LoadQueue.scala 103:51:@5570.10]
  wire  _GEN_600; // @[LoadQueue.scala 104:53:@5571.10]
  wire  _GEN_601; // @[LoadQueue.scala 101:102:@5561.8]
  wire  _GEN_602; // @[LoadQueue.scala 99:27:@5554.6]
  wire  _GEN_603; // @[LoadQueue.scala 95:34:@5539.4]
  wire [4:0] _T_2306; // @[util.scala 10:8:@5582.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@5583.6]
  wire [4:0] _T_2307; // @[util.scala 10:14:@5583.6]
  wire  _T_2308; // @[LoadQueue.scala 97:56:@5584.6]
  wire  _T_2309; // @[LoadQueue.scala 96:50:@5585.6]
  wire  _T_2311; // @[LoadQueue.scala 96:34:@5586.6]
  wire  _T_2313; // @[LoadQueue.scala 101:36:@5594.8]
  wire  _T_2314; // @[LoadQueue.scala 101:86:@5595.8]
  wire  _T_2315; // @[LoadQueue.scala 101:61:@5596.8]
  wire  _T_2318; // @[LoadQueue.scala 103:69:@5602.10]
  wire  _T_2319; // @[LoadQueue.scala 104:31:@5603.10]
  wire  _T_2320; // @[LoadQueue.scala 103:94:@5604.10]
  wire  _T_2322; // @[LoadQueue.scala 103:54:@5605.10]
  wire  _T_2323; // @[LoadQueue.scala 103:51:@5606.10]
  wire  _GEN_620; // @[LoadQueue.scala 104:53:@5607.10]
  wire  _GEN_621; // @[LoadQueue.scala 101:102:@5597.8]
  wire  _GEN_622; // @[LoadQueue.scala 99:27:@5590.6]
  wire  _GEN_623; // @[LoadQueue.scala 95:34:@5575.4]
  wire [4:0] _T_2336; // @[util.scala 10:8:@5618.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@5619.6]
  wire [4:0] _T_2337; // @[util.scala 10:14:@5619.6]
  wire  _T_2338; // @[LoadQueue.scala 97:56:@5620.6]
  wire  _T_2339; // @[LoadQueue.scala 96:50:@5621.6]
  wire  _T_2341; // @[LoadQueue.scala 96:34:@5622.6]
  wire  _T_2343; // @[LoadQueue.scala 101:36:@5630.8]
  wire  _T_2344; // @[LoadQueue.scala 101:86:@5631.8]
  wire  _T_2345; // @[LoadQueue.scala 101:61:@5632.8]
  wire  _T_2348; // @[LoadQueue.scala 103:69:@5638.10]
  wire  _T_2349; // @[LoadQueue.scala 104:31:@5639.10]
  wire  _T_2350; // @[LoadQueue.scala 103:94:@5640.10]
  wire  _T_2352; // @[LoadQueue.scala 103:54:@5641.10]
  wire  _T_2353; // @[LoadQueue.scala 103:51:@5642.10]
  wire  _GEN_640; // @[LoadQueue.scala 104:53:@5643.10]
  wire  _GEN_641; // @[LoadQueue.scala 101:102:@5633.8]
  wire  _GEN_642; // @[LoadQueue.scala 99:27:@5626.6]
  wire  _GEN_643; // @[LoadQueue.scala 95:34:@5611.4]
  wire [4:0] _T_2366; // @[util.scala 10:8:@5654.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@5655.6]
  wire [4:0] _T_2367; // @[util.scala 10:14:@5655.6]
  wire  _T_2368; // @[LoadQueue.scala 97:56:@5656.6]
  wire  _T_2369; // @[LoadQueue.scala 96:50:@5657.6]
  wire  _T_2371; // @[LoadQueue.scala 96:34:@5658.6]
  wire  _T_2373; // @[LoadQueue.scala 101:36:@5666.8]
  wire  _T_2374; // @[LoadQueue.scala 101:86:@5667.8]
  wire  _T_2375; // @[LoadQueue.scala 101:61:@5668.8]
  wire  _T_2378; // @[LoadQueue.scala 103:69:@5674.10]
  wire  _T_2379; // @[LoadQueue.scala 104:31:@5675.10]
  wire  _T_2380; // @[LoadQueue.scala 103:94:@5676.10]
  wire  _T_2382; // @[LoadQueue.scala 103:54:@5677.10]
  wire  _T_2383; // @[LoadQueue.scala 103:51:@5678.10]
  wire  _GEN_660; // @[LoadQueue.scala 104:53:@5679.10]
  wire  _GEN_661; // @[LoadQueue.scala 101:102:@5669.8]
  wire  _GEN_662; // @[LoadQueue.scala 99:27:@5662.6]
  wire  _GEN_663; // @[LoadQueue.scala 95:34:@5647.4]
  wire [4:0] _T_2396; // @[util.scala 10:8:@5690.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@5691.6]
  wire [4:0] _T_2397; // @[util.scala 10:14:@5691.6]
  wire  _T_2398; // @[LoadQueue.scala 97:56:@5692.6]
  wire  _T_2399; // @[LoadQueue.scala 96:50:@5693.6]
  wire  _T_2401; // @[LoadQueue.scala 96:34:@5694.6]
  wire  _T_2403; // @[LoadQueue.scala 101:36:@5702.8]
  wire  _T_2404; // @[LoadQueue.scala 101:86:@5703.8]
  wire  _T_2405; // @[LoadQueue.scala 101:61:@5704.8]
  wire  _T_2408; // @[LoadQueue.scala 103:69:@5710.10]
  wire  _T_2409; // @[LoadQueue.scala 104:31:@5711.10]
  wire  _T_2410; // @[LoadQueue.scala 103:94:@5712.10]
  wire  _T_2412; // @[LoadQueue.scala 103:54:@5713.10]
  wire  _T_2413; // @[LoadQueue.scala 103:51:@5714.10]
  wire  _GEN_680; // @[LoadQueue.scala 104:53:@5715.10]
  wire  _GEN_681; // @[LoadQueue.scala 101:102:@5705.8]
  wire  _GEN_682; // @[LoadQueue.scala 99:27:@5698.6]
  wire  _GEN_683; // @[LoadQueue.scala 95:34:@5683.4]
  wire [4:0] _T_2426; // @[util.scala 10:8:@5726.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@5727.6]
  wire [4:0] _T_2427; // @[util.scala 10:14:@5727.6]
  wire  _T_2428; // @[LoadQueue.scala 97:56:@5728.6]
  wire  _T_2429; // @[LoadQueue.scala 96:50:@5729.6]
  wire  _T_2431; // @[LoadQueue.scala 96:34:@5730.6]
  wire  _T_2433; // @[LoadQueue.scala 101:36:@5738.8]
  wire  _T_2434; // @[LoadQueue.scala 101:86:@5739.8]
  wire  _T_2435; // @[LoadQueue.scala 101:61:@5740.8]
  wire  _T_2438; // @[LoadQueue.scala 103:69:@5746.10]
  wire  _T_2439; // @[LoadQueue.scala 104:31:@5747.10]
  wire  _T_2440; // @[LoadQueue.scala 103:94:@5748.10]
  wire  _T_2442; // @[LoadQueue.scala 103:54:@5749.10]
  wire  _T_2443; // @[LoadQueue.scala 103:51:@5750.10]
  wire  _GEN_700; // @[LoadQueue.scala 104:53:@5751.10]
  wire  _GEN_701; // @[LoadQueue.scala 101:102:@5741.8]
  wire  _GEN_702; // @[LoadQueue.scala 99:27:@5734.6]
  wire  _GEN_703; // @[LoadQueue.scala 95:34:@5719.4]
  wire [4:0] _T_2456; // @[util.scala 10:8:@5762.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@5763.6]
  wire [4:0] _T_2457; // @[util.scala 10:14:@5763.6]
  wire  _T_2458; // @[LoadQueue.scala 97:56:@5764.6]
  wire  _T_2459; // @[LoadQueue.scala 96:50:@5765.6]
  wire  _T_2461; // @[LoadQueue.scala 96:34:@5766.6]
  wire  _T_2463; // @[LoadQueue.scala 101:36:@5774.8]
  wire  _T_2464; // @[LoadQueue.scala 101:86:@5775.8]
  wire  _T_2465; // @[LoadQueue.scala 101:61:@5776.8]
  wire  _T_2468; // @[LoadQueue.scala 103:69:@5782.10]
  wire  _T_2469; // @[LoadQueue.scala 104:31:@5783.10]
  wire  _T_2470; // @[LoadQueue.scala 103:94:@5784.10]
  wire  _T_2472; // @[LoadQueue.scala 103:54:@5785.10]
  wire  _T_2473; // @[LoadQueue.scala 103:51:@5786.10]
  wire  _GEN_720; // @[LoadQueue.scala 104:53:@5787.10]
  wire  _GEN_721; // @[LoadQueue.scala 101:102:@5777.8]
  wire  _GEN_722; // @[LoadQueue.scala 99:27:@5770.6]
  wire  _GEN_723; // @[LoadQueue.scala 95:34:@5755.4]
  wire [4:0] _T_2486; // @[util.scala 10:8:@5798.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@5799.6]
  wire [4:0] _T_2487; // @[util.scala 10:14:@5799.6]
  wire  _T_2488; // @[LoadQueue.scala 97:56:@5800.6]
  wire  _T_2489; // @[LoadQueue.scala 96:50:@5801.6]
  wire  _T_2491; // @[LoadQueue.scala 96:34:@5802.6]
  wire  _T_2493; // @[LoadQueue.scala 101:36:@5810.8]
  wire  _T_2494; // @[LoadQueue.scala 101:86:@5811.8]
  wire  _T_2495; // @[LoadQueue.scala 101:61:@5812.8]
  wire  _T_2498; // @[LoadQueue.scala 103:69:@5818.10]
  wire  _T_2499; // @[LoadQueue.scala 104:31:@5819.10]
  wire  _T_2500; // @[LoadQueue.scala 103:94:@5820.10]
  wire  _T_2502; // @[LoadQueue.scala 103:54:@5821.10]
  wire  _T_2503; // @[LoadQueue.scala 103:51:@5822.10]
  wire  _GEN_740; // @[LoadQueue.scala 104:53:@5823.10]
  wire  _GEN_741; // @[LoadQueue.scala 101:102:@5813.8]
  wire  _GEN_742; // @[LoadQueue.scala 99:27:@5806.6]
  wire  _GEN_743; // @[LoadQueue.scala 95:34:@5791.4]
  wire [4:0] _T_2516; // @[util.scala 10:8:@5834.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@5835.6]
  wire [4:0] _T_2517; // @[util.scala 10:14:@5835.6]
  wire  _T_2518; // @[LoadQueue.scala 97:56:@5836.6]
  wire  _T_2519; // @[LoadQueue.scala 96:50:@5837.6]
  wire  _T_2521; // @[LoadQueue.scala 96:34:@5838.6]
  wire  _T_2523; // @[LoadQueue.scala 101:36:@5846.8]
  wire  _T_2524; // @[LoadQueue.scala 101:86:@5847.8]
  wire  _T_2525; // @[LoadQueue.scala 101:61:@5848.8]
  wire  _T_2528; // @[LoadQueue.scala 103:69:@5854.10]
  wire  _T_2529; // @[LoadQueue.scala 104:31:@5855.10]
  wire  _T_2530; // @[LoadQueue.scala 103:94:@5856.10]
  wire  _T_2532; // @[LoadQueue.scala 103:54:@5857.10]
  wire  _T_2533; // @[LoadQueue.scala 103:51:@5858.10]
  wire  _GEN_760; // @[LoadQueue.scala 104:53:@5859.10]
  wire  _GEN_761; // @[LoadQueue.scala 101:102:@5849.8]
  wire  _GEN_762; // @[LoadQueue.scala 99:27:@5842.6]
  wire  _GEN_763; // @[LoadQueue.scala 95:34:@5827.4]
  wire [4:0] _T_2546; // @[util.scala 10:8:@5870.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@5871.6]
  wire [4:0] _T_2547; // @[util.scala 10:14:@5871.6]
  wire  _T_2548; // @[LoadQueue.scala 97:56:@5872.6]
  wire  _T_2549; // @[LoadQueue.scala 96:50:@5873.6]
  wire  _T_2551; // @[LoadQueue.scala 96:34:@5874.6]
  wire  _T_2553; // @[LoadQueue.scala 101:36:@5882.8]
  wire  _T_2554; // @[LoadQueue.scala 101:86:@5883.8]
  wire  _T_2555; // @[LoadQueue.scala 101:61:@5884.8]
  wire  _T_2558; // @[LoadQueue.scala 103:69:@5890.10]
  wire  _T_2559; // @[LoadQueue.scala 104:31:@5891.10]
  wire  _T_2560; // @[LoadQueue.scala 103:94:@5892.10]
  wire  _T_2562; // @[LoadQueue.scala 103:54:@5893.10]
  wire  _T_2563; // @[LoadQueue.scala 103:51:@5894.10]
  wire  _GEN_780; // @[LoadQueue.scala 104:53:@5895.10]
  wire  _GEN_781; // @[LoadQueue.scala 101:102:@5885.8]
  wire  _GEN_782; // @[LoadQueue.scala 99:27:@5878.6]
  wire  _GEN_783; // @[LoadQueue.scala 95:34:@5863.4]
  wire [4:0] _T_2576; // @[util.scala 10:8:@5906.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@5907.6]
  wire [4:0] _T_2577; // @[util.scala 10:14:@5907.6]
  wire  _T_2578; // @[LoadQueue.scala 97:56:@5908.6]
  wire  _T_2579; // @[LoadQueue.scala 96:50:@5909.6]
  wire  _T_2581; // @[LoadQueue.scala 96:34:@5910.6]
  wire  _T_2583; // @[LoadQueue.scala 101:36:@5918.8]
  wire  _T_2584; // @[LoadQueue.scala 101:86:@5919.8]
  wire  _T_2585; // @[LoadQueue.scala 101:61:@5920.8]
  wire  _T_2588; // @[LoadQueue.scala 103:69:@5926.10]
  wire  _T_2589; // @[LoadQueue.scala 104:31:@5927.10]
  wire  _T_2590; // @[LoadQueue.scala 103:94:@5928.10]
  wire  _T_2592; // @[LoadQueue.scala 103:54:@5929.10]
  wire  _T_2593; // @[LoadQueue.scala 103:51:@5930.10]
  wire  _GEN_800; // @[LoadQueue.scala 104:53:@5931.10]
  wire  _GEN_801; // @[LoadQueue.scala 101:102:@5921.8]
  wire  _GEN_802; // @[LoadQueue.scala 99:27:@5914.6]
  wire  _GEN_803; // @[LoadQueue.scala 95:34:@5899.4]
  wire [4:0] _T_2606; // @[util.scala 10:8:@5942.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@5943.6]
  wire [4:0] _T_2607; // @[util.scala 10:14:@5943.6]
  wire  _T_2608; // @[LoadQueue.scala 97:56:@5944.6]
  wire  _T_2609; // @[LoadQueue.scala 96:50:@5945.6]
  wire  _T_2611; // @[LoadQueue.scala 96:34:@5946.6]
  wire  _T_2613; // @[LoadQueue.scala 101:36:@5954.8]
  wire  _T_2614; // @[LoadQueue.scala 101:86:@5955.8]
  wire  _T_2615; // @[LoadQueue.scala 101:61:@5956.8]
  wire  _T_2618; // @[LoadQueue.scala 103:69:@5962.10]
  wire  _T_2619; // @[LoadQueue.scala 104:31:@5963.10]
  wire  _T_2620; // @[LoadQueue.scala 103:94:@5964.10]
  wire  _T_2622; // @[LoadQueue.scala 103:54:@5965.10]
  wire  _T_2623; // @[LoadQueue.scala 103:51:@5966.10]
  wire  _GEN_820; // @[LoadQueue.scala 104:53:@5967.10]
  wire  _GEN_821; // @[LoadQueue.scala 101:102:@5957.8]
  wire  _GEN_822; // @[LoadQueue.scala 99:27:@5950.6]
  wire  _GEN_823; // @[LoadQueue.scala 95:34:@5935.4]
  wire [4:0] _T_2636; // @[util.scala 10:8:@5978.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@5979.6]
  wire [4:0] _T_2637; // @[util.scala 10:14:@5979.6]
  wire  _T_2638; // @[LoadQueue.scala 97:56:@5980.6]
  wire  _T_2639; // @[LoadQueue.scala 96:50:@5981.6]
  wire  _T_2641; // @[LoadQueue.scala 96:34:@5982.6]
  wire  _T_2643; // @[LoadQueue.scala 101:36:@5990.8]
  wire  _T_2644; // @[LoadQueue.scala 101:86:@5991.8]
  wire  _T_2645; // @[LoadQueue.scala 101:61:@5992.8]
  wire  _T_2648; // @[LoadQueue.scala 103:69:@5998.10]
  wire  _T_2649; // @[LoadQueue.scala 104:31:@5999.10]
  wire  _T_2650; // @[LoadQueue.scala 103:94:@6000.10]
  wire  _T_2652; // @[LoadQueue.scala 103:54:@6001.10]
  wire  _T_2653; // @[LoadQueue.scala 103:51:@6002.10]
  wire  _GEN_840; // @[LoadQueue.scala 104:53:@6003.10]
  wire  _GEN_841; // @[LoadQueue.scala 101:102:@5993.8]
  wire  _GEN_842; // @[LoadQueue.scala 99:27:@5986.6]
  wire  _GEN_843; // @[LoadQueue.scala 95:34:@5971.4]
  wire [4:0] _T_2666; // @[util.scala 10:8:@6014.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@6015.6]
  wire [4:0] _T_2667; // @[util.scala 10:14:@6015.6]
  wire  _T_2668; // @[LoadQueue.scala 97:56:@6016.6]
  wire  _T_2669; // @[LoadQueue.scala 96:50:@6017.6]
  wire  _T_2671; // @[LoadQueue.scala 96:34:@6018.6]
  wire  _T_2673; // @[LoadQueue.scala 101:36:@6026.8]
  wire  _T_2674; // @[LoadQueue.scala 101:86:@6027.8]
  wire  _T_2675; // @[LoadQueue.scala 101:61:@6028.8]
  wire  _T_2678; // @[LoadQueue.scala 103:69:@6034.10]
  wire  _T_2679; // @[LoadQueue.scala 104:31:@6035.10]
  wire  _T_2680; // @[LoadQueue.scala 103:94:@6036.10]
  wire  _T_2682; // @[LoadQueue.scala 103:54:@6037.10]
  wire  _T_2683; // @[LoadQueue.scala 103:51:@6038.10]
  wire  _GEN_860; // @[LoadQueue.scala 104:53:@6039.10]
  wire  _GEN_861; // @[LoadQueue.scala 101:102:@6029.8]
  wire  _GEN_862; // @[LoadQueue.scala 99:27:@6022.6]
  wire  _GEN_863; // @[LoadQueue.scala 95:34:@6007.4]
  wire [15:0] _T_2687; // @[OneHot.scala 52:12:@6044.4]
  wire  _T_2689; // @[util.scala 60:60:@6046.4]
  wire  _T_2690; // @[util.scala 60:60:@6047.4]
  wire  _T_2691; // @[util.scala 60:60:@6048.4]
  wire  _T_2692; // @[util.scala 60:60:@6049.4]
  wire  _T_2693; // @[util.scala 60:60:@6050.4]
  wire  _T_2694; // @[util.scala 60:60:@6051.4]
  wire  _T_2695; // @[util.scala 60:60:@6052.4]
  wire  _T_2696; // @[util.scala 60:60:@6053.4]
  wire  _T_2697; // @[util.scala 60:60:@6054.4]
  wire  _T_2698; // @[util.scala 60:60:@6055.4]
  wire  _T_2699; // @[util.scala 60:60:@6056.4]
  wire  _T_2700; // @[util.scala 60:60:@6057.4]
  wire  _T_2701; // @[util.scala 60:60:@6058.4]
  wire  _T_2702; // @[util.scala 60:60:@6059.4]
  wire  _T_2703; // @[util.scala 60:60:@6060.4]
  wire  _T_2704; // @[util.scala 60:60:@6061.4]
  wire [255:0] _T_4835; // @[Mux.scala 19:72:@7585.4]
  wire [255:0] _T_4842; // @[Mux.scala 19:72:@7592.4]
  wire [511:0] _T_4843; // @[Mux.scala 19:72:@7593.4]
  wire [511:0] _T_4845; // @[Mux.scala 19:72:@7594.4]
  wire [255:0] _T_4852; // @[Mux.scala 19:72:@7601.4]
  wire [255:0] _T_4859; // @[Mux.scala 19:72:@7608.4]
  wire [511:0] _T_4860; // @[Mux.scala 19:72:@7609.4]
  wire [511:0] _T_4862; // @[Mux.scala 19:72:@7610.4]
  wire [255:0] _T_4869; // @[Mux.scala 19:72:@7617.4]
  wire [255:0] _T_4876; // @[Mux.scala 19:72:@7624.4]
  wire [511:0] _T_4877; // @[Mux.scala 19:72:@7625.4]
  wire [511:0] _T_4879; // @[Mux.scala 19:72:@7626.4]
  wire [255:0] _T_4886; // @[Mux.scala 19:72:@7633.4]
  wire [255:0] _T_4893; // @[Mux.scala 19:72:@7640.4]
  wire [511:0] _T_4894; // @[Mux.scala 19:72:@7641.4]
  wire [511:0] _T_4896; // @[Mux.scala 19:72:@7642.4]
  wire [255:0] _T_4903; // @[Mux.scala 19:72:@7649.4]
  wire [255:0] _T_4910; // @[Mux.scala 19:72:@7656.4]
  wire [511:0] _T_4911; // @[Mux.scala 19:72:@7657.4]
  wire [511:0] _T_4913; // @[Mux.scala 19:72:@7658.4]
  wire [255:0] _T_4920; // @[Mux.scala 19:72:@7665.4]
  wire [255:0] _T_4927; // @[Mux.scala 19:72:@7672.4]
  wire [511:0] _T_4928; // @[Mux.scala 19:72:@7673.4]
  wire [511:0] _T_4930; // @[Mux.scala 19:72:@7674.4]
  wire [255:0] _T_4937; // @[Mux.scala 19:72:@7681.4]
  wire [255:0] _T_4944; // @[Mux.scala 19:72:@7688.4]
  wire [511:0] _T_4945; // @[Mux.scala 19:72:@7689.4]
  wire [511:0] _T_4947; // @[Mux.scala 19:72:@7690.4]
  wire [255:0] _T_4954; // @[Mux.scala 19:72:@7697.4]
  wire [255:0] _T_4961; // @[Mux.scala 19:72:@7704.4]
  wire [511:0] _T_4962; // @[Mux.scala 19:72:@7705.4]
  wire [511:0] _T_4964; // @[Mux.scala 19:72:@7706.4]
  wire [511:0] _T_4979; // @[Mux.scala 19:72:@7721.4]
  wire [511:0] _T_4981; // @[Mux.scala 19:72:@7722.4]
  wire [511:0] _T_4996; // @[Mux.scala 19:72:@7737.4]
  wire [511:0] _T_4998; // @[Mux.scala 19:72:@7738.4]
  wire [511:0] _T_5013; // @[Mux.scala 19:72:@7753.4]
  wire [511:0] _T_5015; // @[Mux.scala 19:72:@7754.4]
  wire [511:0] _T_5030; // @[Mux.scala 19:72:@7769.4]
  wire [511:0] _T_5032; // @[Mux.scala 19:72:@7770.4]
  wire [511:0] _T_5047; // @[Mux.scala 19:72:@7785.4]
  wire [511:0] _T_5049; // @[Mux.scala 19:72:@7786.4]
  wire [511:0] _T_5064; // @[Mux.scala 19:72:@7801.4]
  wire [511:0] _T_5066; // @[Mux.scala 19:72:@7802.4]
  wire [511:0] _T_5081; // @[Mux.scala 19:72:@7817.4]
  wire [511:0] _T_5083; // @[Mux.scala 19:72:@7818.4]
  wire [511:0] _T_5098; // @[Mux.scala 19:72:@7833.4]
  wire [511:0] _T_5100; // @[Mux.scala 19:72:@7834.4]
  wire [511:0] _T_5101; // @[Mux.scala 19:72:@7835.4]
  wire [511:0] _T_5102; // @[Mux.scala 19:72:@7836.4]
  wire [511:0] _T_5103; // @[Mux.scala 19:72:@7837.4]
  wire [511:0] _T_5104; // @[Mux.scala 19:72:@7838.4]
  wire [511:0] _T_5105; // @[Mux.scala 19:72:@7839.4]
  wire [511:0] _T_5106; // @[Mux.scala 19:72:@7840.4]
  wire [511:0] _T_5107; // @[Mux.scala 19:72:@7841.4]
  wire [511:0] _T_5108; // @[Mux.scala 19:72:@7842.4]
  wire [511:0] _T_5109; // @[Mux.scala 19:72:@7843.4]
  wire [511:0] _T_5110; // @[Mux.scala 19:72:@7844.4]
  wire [511:0] _T_5111; // @[Mux.scala 19:72:@7845.4]
  wire [511:0] _T_5112; // @[Mux.scala 19:72:@7846.4]
  wire [511:0] _T_5113; // @[Mux.scala 19:72:@7847.4]
  wire [511:0] _T_5114; // @[Mux.scala 19:72:@7848.4]
  wire [511:0] _T_5115; // @[Mux.scala 19:72:@7849.4]
  wire [7:0] _T_5692; // @[Mux.scala 19:72:@8199.4]
  wire [7:0] _T_5699; // @[Mux.scala 19:72:@8206.4]
  wire [15:0] _T_5700; // @[Mux.scala 19:72:@8207.4]
  wire [15:0] _T_5702; // @[Mux.scala 19:72:@8208.4]
  wire [7:0] _T_5709; // @[Mux.scala 19:72:@8215.4]
  wire [7:0] _T_5716; // @[Mux.scala 19:72:@8222.4]
  wire [15:0] _T_5717; // @[Mux.scala 19:72:@8223.4]
  wire [15:0] _T_5719; // @[Mux.scala 19:72:@8224.4]
  wire [7:0] _T_5726; // @[Mux.scala 19:72:@8231.4]
  wire [7:0] _T_5733; // @[Mux.scala 19:72:@8238.4]
  wire [15:0] _T_5734; // @[Mux.scala 19:72:@8239.4]
  wire [15:0] _T_5736; // @[Mux.scala 19:72:@8240.4]
  wire [7:0] _T_5743; // @[Mux.scala 19:72:@8247.4]
  wire [7:0] _T_5750; // @[Mux.scala 19:72:@8254.4]
  wire [15:0] _T_5751; // @[Mux.scala 19:72:@8255.4]
  wire [15:0] _T_5753; // @[Mux.scala 19:72:@8256.4]
  wire [7:0] _T_5760; // @[Mux.scala 19:72:@8263.4]
  wire [7:0] _T_5767; // @[Mux.scala 19:72:@8270.4]
  wire [15:0] _T_5768; // @[Mux.scala 19:72:@8271.4]
  wire [15:0] _T_5770; // @[Mux.scala 19:72:@8272.4]
  wire [7:0] _T_5777; // @[Mux.scala 19:72:@8279.4]
  wire [7:0] _T_5784; // @[Mux.scala 19:72:@8286.4]
  wire [15:0] _T_5785; // @[Mux.scala 19:72:@8287.4]
  wire [15:0] _T_5787; // @[Mux.scala 19:72:@8288.4]
  wire [7:0] _T_5794; // @[Mux.scala 19:72:@8295.4]
  wire [7:0] _T_5801; // @[Mux.scala 19:72:@8302.4]
  wire [15:0] _T_5802; // @[Mux.scala 19:72:@8303.4]
  wire [15:0] _T_5804; // @[Mux.scala 19:72:@8304.4]
  wire [7:0] _T_5811; // @[Mux.scala 19:72:@8311.4]
  wire [7:0] _T_5818; // @[Mux.scala 19:72:@8318.4]
  wire [15:0] _T_5819; // @[Mux.scala 19:72:@8319.4]
  wire [15:0] _T_5821; // @[Mux.scala 19:72:@8320.4]
  wire [15:0] _T_5836; // @[Mux.scala 19:72:@8335.4]
  wire [15:0] _T_5838; // @[Mux.scala 19:72:@8336.4]
  wire [15:0] _T_5853; // @[Mux.scala 19:72:@8351.4]
  wire [15:0] _T_5855; // @[Mux.scala 19:72:@8352.4]
  wire [15:0] _T_5870; // @[Mux.scala 19:72:@8367.4]
  wire [15:0] _T_5872; // @[Mux.scala 19:72:@8368.4]
  wire [15:0] _T_5887; // @[Mux.scala 19:72:@8383.4]
  wire [15:0] _T_5889; // @[Mux.scala 19:72:@8384.4]
  wire [15:0] _T_5904; // @[Mux.scala 19:72:@8399.4]
  wire [15:0] _T_5906; // @[Mux.scala 19:72:@8400.4]
  wire [15:0] _T_5921; // @[Mux.scala 19:72:@8415.4]
  wire [15:0] _T_5923; // @[Mux.scala 19:72:@8416.4]
  wire [15:0] _T_5938; // @[Mux.scala 19:72:@8431.4]
  wire [15:0] _T_5940; // @[Mux.scala 19:72:@8432.4]
  wire [15:0] _T_5955; // @[Mux.scala 19:72:@8447.4]
  wire [15:0] _T_5957; // @[Mux.scala 19:72:@8448.4]
  wire [15:0] _T_5958; // @[Mux.scala 19:72:@8449.4]
  wire [15:0] _T_5959; // @[Mux.scala 19:72:@8450.4]
  wire [15:0] _T_5960; // @[Mux.scala 19:72:@8451.4]
  wire [15:0] _T_5961; // @[Mux.scala 19:72:@8452.4]
  wire [15:0] _T_5962; // @[Mux.scala 19:72:@8453.4]
  wire [15:0] _T_5963; // @[Mux.scala 19:72:@8454.4]
  wire [15:0] _T_5964; // @[Mux.scala 19:72:@8455.4]
  wire [15:0] _T_5965; // @[Mux.scala 19:72:@8456.4]
  wire [15:0] _T_5966; // @[Mux.scala 19:72:@8457.4]
  wire [15:0] _T_5967; // @[Mux.scala 19:72:@8458.4]
  wire [15:0] _T_5968; // @[Mux.scala 19:72:@8459.4]
  wire [15:0] _T_5969; // @[Mux.scala 19:72:@8460.4]
  wire [15:0] _T_5970; // @[Mux.scala 19:72:@8461.4]
  wire [15:0] _T_5971; // @[Mux.scala 19:72:@8462.4]
  wire [15:0] _T_5972; // @[Mux.scala 19:72:@8463.4]
  wire  _T_6113; // @[LoadQueue.scala 121:105:@8499.4]
  wire  _T_6115; // @[LoadQueue.scala 122:18:@8500.4]
  wire  _T_6117; // @[LoadQueue.scala 122:36:@8501.4]
  wire  _T_6118; // @[LoadQueue.scala 122:27:@8502.4]
  wire  _T_6120; // @[LoadQueue.scala 122:52:@8503.4]
  wire  _T_6122; // @[LoadQueue.scala 122:85:@8504.4]
  wire  _T_6124; // @[LoadQueue.scala 122:103:@8505.4]
  wire  _T_6125; // @[LoadQueue.scala 122:94:@8506.4]
  wire  _T_6127; // @[LoadQueue.scala 122:70:@8507.4]
  wire  _T_6128; // @[LoadQueue.scala 122:67:@8508.4]
  wire  validEntriesInStoreQ_0; // @[LoadQueue.scala 121:91:@8509.4]
  wire  _T_6132; // @[LoadQueue.scala 122:18:@8511.4]
  wire  _T_6134; // @[LoadQueue.scala 122:36:@8512.4]
  wire  _T_6135; // @[LoadQueue.scala 122:27:@8513.4]
  wire  _T_6139; // @[LoadQueue.scala 122:85:@8515.4]
  wire  _T_6141; // @[LoadQueue.scala 122:103:@8516.4]
  wire  _T_6142; // @[LoadQueue.scala 122:94:@8517.4]
  wire  _T_6144; // @[LoadQueue.scala 122:70:@8518.4]
  wire  _T_6145; // @[LoadQueue.scala 122:67:@8519.4]
  wire  validEntriesInStoreQ_1; // @[LoadQueue.scala 121:91:@8520.4]
  wire  _T_6149; // @[LoadQueue.scala 122:18:@8522.4]
  wire  _T_6151; // @[LoadQueue.scala 122:36:@8523.4]
  wire  _T_6152; // @[LoadQueue.scala 122:27:@8524.4]
  wire  _T_6156; // @[LoadQueue.scala 122:85:@8526.4]
  wire  _T_6158; // @[LoadQueue.scala 122:103:@8527.4]
  wire  _T_6159; // @[LoadQueue.scala 122:94:@8528.4]
  wire  _T_6161; // @[LoadQueue.scala 122:70:@8529.4]
  wire  _T_6162; // @[LoadQueue.scala 122:67:@8530.4]
  wire  validEntriesInStoreQ_2; // @[LoadQueue.scala 121:91:@8531.4]
  wire  _T_6166; // @[LoadQueue.scala 122:18:@8533.4]
  wire  _T_6168; // @[LoadQueue.scala 122:36:@8534.4]
  wire  _T_6169; // @[LoadQueue.scala 122:27:@8535.4]
  wire  _T_6173; // @[LoadQueue.scala 122:85:@8537.4]
  wire  _T_6175; // @[LoadQueue.scala 122:103:@8538.4]
  wire  _T_6176; // @[LoadQueue.scala 122:94:@8539.4]
  wire  _T_6178; // @[LoadQueue.scala 122:70:@8540.4]
  wire  _T_6179; // @[LoadQueue.scala 122:67:@8541.4]
  wire  validEntriesInStoreQ_3; // @[LoadQueue.scala 121:91:@8542.4]
  wire  _T_6183; // @[LoadQueue.scala 122:18:@8544.4]
  wire  _T_6185; // @[LoadQueue.scala 122:36:@8545.4]
  wire  _T_6186; // @[LoadQueue.scala 122:27:@8546.4]
  wire  _T_6190; // @[LoadQueue.scala 122:85:@8548.4]
  wire  _T_6192; // @[LoadQueue.scala 122:103:@8549.4]
  wire  _T_6193; // @[LoadQueue.scala 122:94:@8550.4]
  wire  _T_6195; // @[LoadQueue.scala 122:70:@8551.4]
  wire  _T_6196; // @[LoadQueue.scala 122:67:@8552.4]
  wire  validEntriesInStoreQ_4; // @[LoadQueue.scala 121:91:@8553.4]
  wire  _T_6200; // @[LoadQueue.scala 122:18:@8555.4]
  wire  _T_6202; // @[LoadQueue.scala 122:36:@8556.4]
  wire  _T_6203; // @[LoadQueue.scala 122:27:@8557.4]
  wire  _T_6207; // @[LoadQueue.scala 122:85:@8559.4]
  wire  _T_6209; // @[LoadQueue.scala 122:103:@8560.4]
  wire  _T_6210; // @[LoadQueue.scala 122:94:@8561.4]
  wire  _T_6212; // @[LoadQueue.scala 122:70:@8562.4]
  wire  _T_6213; // @[LoadQueue.scala 122:67:@8563.4]
  wire  validEntriesInStoreQ_5; // @[LoadQueue.scala 121:91:@8564.4]
  wire  _T_6217; // @[LoadQueue.scala 122:18:@8566.4]
  wire  _T_6219; // @[LoadQueue.scala 122:36:@8567.4]
  wire  _T_6220; // @[LoadQueue.scala 122:27:@8568.4]
  wire  _T_6224; // @[LoadQueue.scala 122:85:@8570.4]
  wire  _T_6226; // @[LoadQueue.scala 122:103:@8571.4]
  wire  _T_6227; // @[LoadQueue.scala 122:94:@8572.4]
  wire  _T_6229; // @[LoadQueue.scala 122:70:@8573.4]
  wire  _T_6230; // @[LoadQueue.scala 122:67:@8574.4]
  wire  validEntriesInStoreQ_6; // @[LoadQueue.scala 121:91:@8575.4]
  wire  _T_6234; // @[LoadQueue.scala 122:18:@8577.4]
  wire  _T_6236; // @[LoadQueue.scala 122:36:@8578.4]
  wire  _T_6237; // @[LoadQueue.scala 122:27:@8579.4]
  wire  _T_6241; // @[LoadQueue.scala 122:85:@8581.4]
  wire  _T_6243; // @[LoadQueue.scala 122:103:@8582.4]
  wire  _T_6244; // @[LoadQueue.scala 122:94:@8583.4]
  wire  _T_6246; // @[LoadQueue.scala 122:70:@8584.4]
  wire  _T_6247; // @[LoadQueue.scala 122:67:@8585.4]
  wire  validEntriesInStoreQ_7; // @[LoadQueue.scala 121:91:@8586.4]
  wire  _T_6251; // @[LoadQueue.scala 122:18:@8588.4]
  wire  _T_6253; // @[LoadQueue.scala 122:36:@8589.4]
  wire  _T_6254; // @[LoadQueue.scala 122:27:@8590.4]
  wire  _T_6258; // @[LoadQueue.scala 122:85:@8592.4]
  wire  _T_6260; // @[LoadQueue.scala 122:103:@8593.4]
  wire  _T_6261; // @[LoadQueue.scala 122:94:@8594.4]
  wire  _T_6263; // @[LoadQueue.scala 122:70:@8595.4]
  wire  _T_6264; // @[LoadQueue.scala 122:67:@8596.4]
  wire  validEntriesInStoreQ_8; // @[LoadQueue.scala 121:91:@8597.4]
  wire  _T_6268; // @[LoadQueue.scala 122:18:@8599.4]
  wire  _T_6270; // @[LoadQueue.scala 122:36:@8600.4]
  wire  _T_6271; // @[LoadQueue.scala 122:27:@8601.4]
  wire  _T_6275; // @[LoadQueue.scala 122:85:@8603.4]
  wire  _T_6277; // @[LoadQueue.scala 122:103:@8604.4]
  wire  _T_6278; // @[LoadQueue.scala 122:94:@8605.4]
  wire  _T_6280; // @[LoadQueue.scala 122:70:@8606.4]
  wire  _T_6281; // @[LoadQueue.scala 122:67:@8607.4]
  wire  validEntriesInStoreQ_9; // @[LoadQueue.scala 121:91:@8608.4]
  wire  _T_6285; // @[LoadQueue.scala 122:18:@8610.4]
  wire  _T_6287; // @[LoadQueue.scala 122:36:@8611.4]
  wire  _T_6288; // @[LoadQueue.scala 122:27:@8612.4]
  wire  _T_6292; // @[LoadQueue.scala 122:85:@8614.4]
  wire  _T_6294; // @[LoadQueue.scala 122:103:@8615.4]
  wire  _T_6295; // @[LoadQueue.scala 122:94:@8616.4]
  wire  _T_6297; // @[LoadQueue.scala 122:70:@8617.4]
  wire  _T_6298; // @[LoadQueue.scala 122:67:@8618.4]
  wire  validEntriesInStoreQ_10; // @[LoadQueue.scala 121:91:@8619.4]
  wire  _T_6302; // @[LoadQueue.scala 122:18:@8621.4]
  wire  _T_6304; // @[LoadQueue.scala 122:36:@8622.4]
  wire  _T_6305; // @[LoadQueue.scala 122:27:@8623.4]
  wire  _T_6309; // @[LoadQueue.scala 122:85:@8625.4]
  wire  _T_6311; // @[LoadQueue.scala 122:103:@8626.4]
  wire  _T_6312; // @[LoadQueue.scala 122:94:@8627.4]
  wire  _T_6314; // @[LoadQueue.scala 122:70:@8628.4]
  wire  _T_6315; // @[LoadQueue.scala 122:67:@8629.4]
  wire  validEntriesInStoreQ_11; // @[LoadQueue.scala 121:91:@8630.4]
  wire  _T_6319; // @[LoadQueue.scala 122:18:@8632.4]
  wire  _T_6321; // @[LoadQueue.scala 122:36:@8633.4]
  wire  _T_6322; // @[LoadQueue.scala 122:27:@8634.4]
  wire  _T_6326; // @[LoadQueue.scala 122:85:@8636.4]
  wire  _T_6328; // @[LoadQueue.scala 122:103:@8637.4]
  wire  _T_6329; // @[LoadQueue.scala 122:94:@8638.4]
  wire  _T_6331; // @[LoadQueue.scala 122:70:@8639.4]
  wire  _T_6332; // @[LoadQueue.scala 122:67:@8640.4]
  wire  validEntriesInStoreQ_12; // @[LoadQueue.scala 121:91:@8641.4]
  wire  _T_6336; // @[LoadQueue.scala 122:18:@8643.4]
  wire  _T_6338; // @[LoadQueue.scala 122:36:@8644.4]
  wire  _T_6339; // @[LoadQueue.scala 122:27:@8645.4]
  wire  _T_6343; // @[LoadQueue.scala 122:85:@8647.4]
  wire  _T_6345; // @[LoadQueue.scala 122:103:@8648.4]
  wire  _T_6346; // @[LoadQueue.scala 122:94:@8649.4]
  wire  _T_6348; // @[LoadQueue.scala 122:70:@8650.4]
  wire  _T_6349; // @[LoadQueue.scala 122:67:@8651.4]
  wire  validEntriesInStoreQ_13; // @[LoadQueue.scala 121:91:@8652.4]
  wire  _T_6353; // @[LoadQueue.scala 122:18:@8654.4]
  wire  _T_6355; // @[LoadQueue.scala 122:36:@8655.4]
  wire  _T_6356; // @[LoadQueue.scala 122:27:@8656.4]
  wire  _T_6360; // @[LoadQueue.scala 122:85:@8658.4]
  wire  _T_6362; // @[LoadQueue.scala 122:103:@8659.4]
  wire  _T_6363; // @[LoadQueue.scala 122:94:@8660.4]
  wire  _T_6365; // @[LoadQueue.scala 122:70:@8661.4]
  wire  _T_6366; // @[LoadQueue.scala 122:67:@8662.4]
  wire  validEntriesInStoreQ_14; // @[LoadQueue.scala 121:91:@8663.4]
  wire  validEntriesInStoreQ_15; // @[LoadQueue.scala 121:91:@8674.4]
  wire  storesToCheck_0_0; // @[LoadQueue.scala 131:10:@8701.4]
  wire  _T_7654; // @[LoadQueue.scala 131:81:@8704.4]
  wire  _T_7655; // @[LoadQueue.scala 131:72:@8705.4]
  wire  _T_7657; // @[LoadQueue.scala 132:33:@8706.4]
  wire  _T_7660; // @[LoadQueue.scala 132:41:@8708.4]
  wire  _T_7662; // @[LoadQueue.scala 132:9:@8709.4]
  wire  storesToCheck_0_1; // @[LoadQueue.scala 131:10:@8710.4]
  wire  _T_7668; // @[LoadQueue.scala 131:81:@8713.4]
  wire  _T_7669; // @[LoadQueue.scala 131:72:@8714.4]
  wire  _T_7671; // @[LoadQueue.scala 132:33:@8715.4]
  wire  _T_7674; // @[LoadQueue.scala 132:41:@8717.4]
  wire  _T_7676; // @[LoadQueue.scala 132:9:@8718.4]
  wire  storesToCheck_0_2; // @[LoadQueue.scala 131:10:@8719.4]
  wire  _T_7682; // @[LoadQueue.scala 131:81:@8722.4]
  wire  _T_7683; // @[LoadQueue.scala 131:72:@8723.4]
  wire  _T_7685; // @[LoadQueue.scala 132:33:@8724.4]
  wire  _T_7688; // @[LoadQueue.scala 132:41:@8726.4]
  wire  _T_7690; // @[LoadQueue.scala 132:9:@8727.4]
  wire  storesToCheck_0_3; // @[LoadQueue.scala 131:10:@8728.4]
  wire  _T_7696; // @[LoadQueue.scala 131:81:@8731.4]
  wire  _T_7697; // @[LoadQueue.scala 131:72:@8732.4]
  wire  _T_7699; // @[LoadQueue.scala 132:33:@8733.4]
  wire  _T_7702; // @[LoadQueue.scala 132:41:@8735.4]
  wire  _T_7704; // @[LoadQueue.scala 132:9:@8736.4]
  wire  storesToCheck_0_4; // @[LoadQueue.scala 131:10:@8737.4]
  wire  _T_7710; // @[LoadQueue.scala 131:81:@8740.4]
  wire  _T_7711; // @[LoadQueue.scala 131:72:@8741.4]
  wire  _T_7713; // @[LoadQueue.scala 132:33:@8742.4]
  wire  _T_7716; // @[LoadQueue.scala 132:41:@8744.4]
  wire  _T_7718; // @[LoadQueue.scala 132:9:@8745.4]
  wire  storesToCheck_0_5; // @[LoadQueue.scala 131:10:@8746.4]
  wire  _T_7724; // @[LoadQueue.scala 131:81:@8749.4]
  wire  _T_7725; // @[LoadQueue.scala 131:72:@8750.4]
  wire  _T_7727; // @[LoadQueue.scala 132:33:@8751.4]
  wire  _T_7730; // @[LoadQueue.scala 132:41:@8753.4]
  wire  _T_7732; // @[LoadQueue.scala 132:9:@8754.4]
  wire  storesToCheck_0_6; // @[LoadQueue.scala 131:10:@8755.4]
  wire  _T_7738; // @[LoadQueue.scala 131:81:@8758.4]
  wire  _T_7739; // @[LoadQueue.scala 131:72:@8759.4]
  wire  _T_7741; // @[LoadQueue.scala 132:33:@8760.4]
  wire  _T_7744; // @[LoadQueue.scala 132:41:@8762.4]
  wire  _T_7746; // @[LoadQueue.scala 132:9:@8763.4]
  wire  storesToCheck_0_7; // @[LoadQueue.scala 131:10:@8764.4]
  wire  _T_7752; // @[LoadQueue.scala 131:81:@8767.4]
  wire  _T_7753; // @[LoadQueue.scala 131:72:@8768.4]
  wire  _T_7755; // @[LoadQueue.scala 132:33:@8769.4]
  wire  _T_7758; // @[LoadQueue.scala 132:41:@8771.4]
  wire  _T_7760; // @[LoadQueue.scala 132:9:@8772.4]
  wire  storesToCheck_0_8; // @[LoadQueue.scala 131:10:@8773.4]
  wire  _T_7766; // @[LoadQueue.scala 131:81:@8776.4]
  wire  _T_7767; // @[LoadQueue.scala 131:72:@8777.4]
  wire  _T_7769; // @[LoadQueue.scala 132:33:@8778.4]
  wire  _T_7772; // @[LoadQueue.scala 132:41:@8780.4]
  wire  _T_7774; // @[LoadQueue.scala 132:9:@8781.4]
  wire  storesToCheck_0_9; // @[LoadQueue.scala 131:10:@8782.4]
  wire  _T_7780; // @[LoadQueue.scala 131:81:@8785.4]
  wire  _T_7781; // @[LoadQueue.scala 131:72:@8786.4]
  wire  _T_7783; // @[LoadQueue.scala 132:33:@8787.4]
  wire  _T_7786; // @[LoadQueue.scala 132:41:@8789.4]
  wire  _T_7788; // @[LoadQueue.scala 132:9:@8790.4]
  wire  storesToCheck_0_10; // @[LoadQueue.scala 131:10:@8791.4]
  wire  _T_7794; // @[LoadQueue.scala 131:81:@8794.4]
  wire  _T_7795; // @[LoadQueue.scala 131:72:@8795.4]
  wire  _T_7797; // @[LoadQueue.scala 132:33:@8796.4]
  wire  _T_7800; // @[LoadQueue.scala 132:41:@8798.4]
  wire  _T_7802; // @[LoadQueue.scala 132:9:@8799.4]
  wire  storesToCheck_0_11; // @[LoadQueue.scala 131:10:@8800.4]
  wire  _T_7808; // @[LoadQueue.scala 131:81:@8803.4]
  wire  _T_7809; // @[LoadQueue.scala 131:72:@8804.4]
  wire  _T_7811; // @[LoadQueue.scala 132:33:@8805.4]
  wire  _T_7814; // @[LoadQueue.scala 132:41:@8807.4]
  wire  _T_7816; // @[LoadQueue.scala 132:9:@8808.4]
  wire  storesToCheck_0_12; // @[LoadQueue.scala 131:10:@8809.4]
  wire  _T_7822; // @[LoadQueue.scala 131:81:@8812.4]
  wire  _T_7823; // @[LoadQueue.scala 131:72:@8813.4]
  wire  _T_7825; // @[LoadQueue.scala 132:33:@8814.4]
  wire  _T_7828; // @[LoadQueue.scala 132:41:@8816.4]
  wire  _T_7830; // @[LoadQueue.scala 132:9:@8817.4]
  wire  storesToCheck_0_13; // @[LoadQueue.scala 131:10:@8818.4]
  wire  _T_7836; // @[LoadQueue.scala 131:81:@8821.4]
  wire  _T_7837; // @[LoadQueue.scala 131:72:@8822.4]
  wire  _T_7839; // @[LoadQueue.scala 132:33:@8823.4]
  wire  _T_7842; // @[LoadQueue.scala 132:41:@8825.4]
  wire  _T_7844; // @[LoadQueue.scala 132:9:@8826.4]
  wire  storesToCheck_0_14; // @[LoadQueue.scala 131:10:@8827.4]
  wire  _T_7850; // @[LoadQueue.scala 131:81:@8830.4]
  wire  storesToCheck_0_15; // @[LoadQueue.scala 131:10:@8836.4]
  wire  storesToCheck_1_0; // @[LoadQueue.scala 131:10:@8878.4]
  wire  _T_7900; // @[LoadQueue.scala 131:81:@8881.4]
  wire  _T_7901; // @[LoadQueue.scala 131:72:@8882.4]
  wire  _T_7903; // @[LoadQueue.scala 132:33:@8883.4]
  wire  _T_7906; // @[LoadQueue.scala 132:41:@8885.4]
  wire  _T_7908; // @[LoadQueue.scala 132:9:@8886.4]
  wire  storesToCheck_1_1; // @[LoadQueue.scala 131:10:@8887.4]
  wire  _T_7914; // @[LoadQueue.scala 131:81:@8890.4]
  wire  _T_7915; // @[LoadQueue.scala 131:72:@8891.4]
  wire  _T_7917; // @[LoadQueue.scala 132:33:@8892.4]
  wire  _T_7920; // @[LoadQueue.scala 132:41:@8894.4]
  wire  _T_7922; // @[LoadQueue.scala 132:9:@8895.4]
  wire  storesToCheck_1_2; // @[LoadQueue.scala 131:10:@8896.4]
  wire  _T_7928; // @[LoadQueue.scala 131:81:@8899.4]
  wire  _T_7929; // @[LoadQueue.scala 131:72:@8900.4]
  wire  _T_7931; // @[LoadQueue.scala 132:33:@8901.4]
  wire  _T_7934; // @[LoadQueue.scala 132:41:@8903.4]
  wire  _T_7936; // @[LoadQueue.scala 132:9:@8904.4]
  wire  storesToCheck_1_3; // @[LoadQueue.scala 131:10:@8905.4]
  wire  _T_7942; // @[LoadQueue.scala 131:81:@8908.4]
  wire  _T_7943; // @[LoadQueue.scala 131:72:@8909.4]
  wire  _T_7945; // @[LoadQueue.scala 132:33:@8910.4]
  wire  _T_7948; // @[LoadQueue.scala 132:41:@8912.4]
  wire  _T_7950; // @[LoadQueue.scala 132:9:@8913.4]
  wire  storesToCheck_1_4; // @[LoadQueue.scala 131:10:@8914.4]
  wire  _T_7956; // @[LoadQueue.scala 131:81:@8917.4]
  wire  _T_7957; // @[LoadQueue.scala 131:72:@8918.4]
  wire  _T_7959; // @[LoadQueue.scala 132:33:@8919.4]
  wire  _T_7962; // @[LoadQueue.scala 132:41:@8921.4]
  wire  _T_7964; // @[LoadQueue.scala 132:9:@8922.4]
  wire  storesToCheck_1_5; // @[LoadQueue.scala 131:10:@8923.4]
  wire  _T_7970; // @[LoadQueue.scala 131:81:@8926.4]
  wire  _T_7971; // @[LoadQueue.scala 131:72:@8927.4]
  wire  _T_7973; // @[LoadQueue.scala 132:33:@8928.4]
  wire  _T_7976; // @[LoadQueue.scala 132:41:@8930.4]
  wire  _T_7978; // @[LoadQueue.scala 132:9:@8931.4]
  wire  storesToCheck_1_6; // @[LoadQueue.scala 131:10:@8932.4]
  wire  _T_7984; // @[LoadQueue.scala 131:81:@8935.4]
  wire  _T_7985; // @[LoadQueue.scala 131:72:@8936.4]
  wire  _T_7987; // @[LoadQueue.scala 132:33:@8937.4]
  wire  _T_7990; // @[LoadQueue.scala 132:41:@8939.4]
  wire  _T_7992; // @[LoadQueue.scala 132:9:@8940.4]
  wire  storesToCheck_1_7; // @[LoadQueue.scala 131:10:@8941.4]
  wire  _T_7998; // @[LoadQueue.scala 131:81:@8944.4]
  wire  _T_7999; // @[LoadQueue.scala 131:72:@8945.4]
  wire  _T_8001; // @[LoadQueue.scala 132:33:@8946.4]
  wire  _T_8004; // @[LoadQueue.scala 132:41:@8948.4]
  wire  _T_8006; // @[LoadQueue.scala 132:9:@8949.4]
  wire  storesToCheck_1_8; // @[LoadQueue.scala 131:10:@8950.4]
  wire  _T_8012; // @[LoadQueue.scala 131:81:@8953.4]
  wire  _T_8013; // @[LoadQueue.scala 131:72:@8954.4]
  wire  _T_8015; // @[LoadQueue.scala 132:33:@8955.4]
  wire  _T_8018; // @[LoadQueue.scala 132:41:@8957.4]
  wire  _T_8020; // @[LoadQueue.scala 132:9:@8958.4]
  wire  storesToCheck_1_9; // @[LoadQueue.scala 131:10:@8959.4]
  wire  _T_8026; // @[LoadQueue.scala 131:81:@8962.4]
  wire  _T_8027; // @[LoadQueue.scala 131:72:@8963.4]
  wire  _T_8029; // @[LoadQueue.scala 132:33:@8964.4]
  wire  _T_8032; // @[LoadQueue.scala 132:41:@8966.4]
  wire  _T_8034; // @[LoadQueue.scala 132:9:@8967.4]
  wire  storesToCheck_1_10; // @[LoadQueue.scala 131:10:@8968.4]
  wire  _T_8040; // @[LoadQueue.scala 131:81:@8971.4]
  wire  _T_8041; // @[LoadQueue.scala 131:72:@8972.4]
  wire  _T_8043; // @[LoadQueue.scala 132:33:@8973.4]
  wire  _T_8046; // @[LoadQueue.scala 132:41:@8975.4]
  wire  _T_8048; // @[LoadQueue.scala 132:9:@8976.4]
  wire  storesToCheck_1_11; // @[LoadQueue.scala 131:10:@8977.4]
  wire  _T_8054; // @[LoadQueue.scala 131:81:@8980.4]
  wire  _T_8055; // @[LoadQueue.scala 131:72:@8981.4]
  wire  _T_8057; // @[LoadQueue.scala 132:33:@8982.4]
  wire  _T_8060; // @[LoadQueue.scala 132:41:@8984.4]
  wire  _T_8062; // @[LoadQueue.scala 132:9:@8985.4]
  wire  storesToCheck_1_12; // @[LoadQueue.scala 131:10:@8986.4]
  wire  _T_8068; // @[LoadQueue.scala 131:81:@8989.4]
  wire  _T_8069; // @[LoadQueue.scala 131:72:@8990.4]
  wire  _T_8071; // @[LoadQueue.scala 132:33:@8991.4]
  wire  _T_8074; // @[LoadQueue.scala 132:41:@8993.4]
  wire  _T_8076; // @[LoadQueue.scala 132:9:@8994.4]
  wire  storesToCheck_1_13; // @[LoadQueue.scala 131:10:@8995.4]
  wire  _T_8082; // @[LoadQueue.scala 131:81:@8998.4]
  wire  _T_8083; // @[LoadQueue.scala 131:72:@8999.4]
  wire  _T_8085; // @[LoadQueue.scala 132:33:@9000.4]
  wire  _T_8088; // @[LoadQueue.scala 132:41:@9002.4]
  wire  _T_8090; // @[LoadQueue.scala 132:9:@9003.4]
  wire  storesToCheck_1_14; // @[LoadQueue.scala 131:10:@9004.4]
  wire  _T_8096; // @[LoadQueue.scala 131:81:@9007.4]
  wire  storesToCheck_1_15; // @[LoadQueue.scala 131:10:@9013.4]
  wire  storesToCheck_2_0; // @[LoadQueue.scala 131:10:@9055.4]
  wire  _T_8146; // @[LoadQueue.scala 131:81:@9058.4]
  wire  _T_8147; // @[LoadQueue.scala 131:72:@9059.4]
  wire  _T_8149; // @[LoadQueue.scala 132:33:@9060.4]
  wire  _T_8152; // @[LoadQueue.scala 132:41:@9062.4]
  wire  _T_8154; // @[LoadQueue.scala 132:9:@9063.4]
  wire  storesToCheck_2_1; // @[LoadQueue.scala 131:10:@9064.4]
  wire  _T_8160; // @[LoadQueue.scala 131:81:@9067.4]
  wire  _T_8161; // @[LoadQueue.scala 131:72:@9068.4]
  wire  _T_8163; // @[LoadQueue.scala 132:33:@9069.4]
  wire  _T_8166; // @[LoadQueue.scala 132:41:@9071.4]
  wire  _T_8168; // @[LoadQueue.scala 132:9:@9072.4]
  wire  storesToCheck_2_2; // @[LoadQueue.scala 131:10:@9073.4]
  wire  _T_8174; // @[LoadQueue.scala 131:81:@9076.4]
  wire  _T_8175; // @[LoadQueue.scala 131:72:@9077.4]
  wire  _T_8177; // @[LoadQueue.scala 132:33:@9078.4]
  wire  _T_8180; // @[LoadQueue.scala 132:41:@9080.4]
  wire  _T_8182; // @[LoadQueue.scala 132:9:@9081.4]
  wire  storesToCheck_2_3; // @[LoadQueue.scala 131:10:@9082.4]
  wire  _T_8188; // @[LoadQueue.scala 131:81:@9085.4]
  wire  _T_8189; // @[LoadQueue.scala 131:72:@9086.4]
  wire  _T_8191; // @[LoadQueue.scala 132:33:@9087.4]
  wire  _T_8194; // @[LoadQueue.scala 132:41:@9089.4]
  wire  _T_8196; // @[LoadQueue.scala 132:9:@9090.4]
  wire  storesToCheck_2_4; // @[LoadQueue.scala 131:10:@9091.4]
  wire  _T_8202; // @[LoadQueue.scala 131:81:@9094.4]
  wire  _T_8203; // @[LoadQueue.scala 131:72:@9095.4]
  wire  _T_8205; // @[LoadQueue.scala 132:33:@9096.4]
  wire  _T_8208; // @[LoadQueue.scala 132:41:@9098.4]
  wire  _T_8210; // @[LoadQueue.scala 132:9:@9099.4]
  wire  storesToCheck_2_5; // @[LoadQueue.scala 131:10:@9100.4]
  wire  _T_8216; // @[LoadQueue.scala 131:81:@9103.4]
  wire  _T_8217; // @[LoadQueue.scala 131:72:@9104.4]
  wire  _T_8219; // @[LoadQueue.scala 132:33:@9105.4]
  wire  _T_8222; // @[LoadQueue.scala 132:41:@9107.4]
  wire  _T_8224; // @[LoadQueue.scala 132:9:@9108.4]
  wire  storesToCheck_2_6; // @[LoadQueue.scala 131:10:@9109.4]
  wire  _T_8230; // @[LoadQueue.scala 131:81:@9112.4]
  wire  _T_8231; // @[LoadQueue.scala 131:72:@9113.4]
  wire  _T_8233; // @[LoadQueue.scala 132:33:@9114.4]
  wire  _T_8236; // @[LoadQueue.scala 132:41:@9116.4]
  wire  _T_8238; // @[LoadQueue.scala 132:9:@9117.4]
  wire  storesToCheck_2_7; // @[LoadQueue.scala 131:10:@9118.4]
  wire  _T_8244; // @[LoadQueue.scala 131:81:@9121.4]
  wire  _T_8245; // @[LoadQueue.scala 131:72:@9122.4]
  wire  _T_8247; // @[LoadQueue.scala 132:33:@9123.4]
  wire  _T_8250; // @[LoadQueue.scala 132:41:@9125.4]
  wire  _T_8252; // @[LoadQueue.scala 132:9:@9126.4]
  wire  storesToCheck_2_8; // @[LoadQueue.scala 131:10:@9127.4]
  wire  _T_8258; // @[LoadQueue.scala 131:81:@9130.4]
  wire  _T_8259; // @[LoadQueue.scala 131:72:@9131.4]
  wire  _T_8261; // @[LoadQueue.scala 132:33:@9132.4]
  wire  _T_8264; // @[LoadQueue.scala 132:41:@9134.4]
  wire  _T_8266; // @[LoadQueue.scala 132:9:@9135.4]
  wire  storesToCheck_2_9; // @[LoadQueue.scala 131:10:@9136.4]
  wire  _T_8272; // @[LoadQueue.scala 131:81:@9139.4]
  wire  _T_8273; // @[LoadQueue.scala 131:72:@9140.4]
  wire  _T_8275; // @[LoadQueue.scala 132:33:@9141.4]
  wire  _T_8278; // @[LoadQueue.scala 132:41:@9143.4]
  wire  _T_8280; // @[LoadQueue.scala 132:9:@9144.4]
  wire  storesToCheck_2_10; // @[LoadQueue.scala 131:10:@9145.4]
  wire  _T_8286; // @[LoadQueue.scala 131:81:@9148.4]
  wire  _T_8287; // @[LoadQueue.scala 131:72:@9149.4]
  wire  _T_8289; // @[LoadQueue.scala 132:33:@9150.4]
  wire  _T_8292; // @[LoadQueue.scala 132:41:@9152.4]
  wire  _T_8294; // @[LoadQueue.scala 132:9:@9153.4]
  wire  storesToCheck_2_11; // @[LoadQueue.scala 131:10:@9154.4]
  wire  _T_8300; // @[LoadQueue.scala 131:81:@9157.4]
  wire  _T_8301; // @[LoadQueue.scala 131:72:@9158.4]
  wire  _T_8303; // @[LoadQueue.scala 132:33:@9159.4]
  wire  _T_8306; // @[LoadQueue.scala 132:41:@9161.4]
  wire  _T_8308; // @[LoadQueue.scala 132:9:@9162.4]
  wire  storesToCheck_2_12; // @[LoadQueue.scala 131:10:@9163.4]
  wire  _T_8314; // @[LoadQueue.scala 131:81:@9166.4]
  wire  _T_8315; // @[LoadQueue.scala 131:72:@9167.4]
  wire  _T_8317; // @[LoadQueue.scala 132:33:@9168.4]
  wire  _T_8320; // @[LoadQueue.scala 132:41:@9170.4]
  wire  _T_8322; // @[LoadQueue.scala 132:9:@9171.4]
  wire  storesToCheck_2_13; // @[LoadQueue.scala 131:10:@9172.4]
  wire  _T_8328; // @[LoadQueue.scala 131:81:@9175.4]
  wire  _T_8329; // @[LoadQueue.scala 131:72:@9176.4]
  wire  _T_8331; // @[LoadQueue.scala 132:33:@9177.4]
  wire  _T_8334; // @[LoadQueue.scala 132:41:@9179.4]
  wire  _T_8336; // @[LoadQueue.scala 132:9:@9180.4]
  wire  storesToCheck_2_14; // @[LoadQueue.scala 131:10:@9181.4]
  wire  _T_8342; // @[LoadQueue.scala 131:81:@9184.4]
  wire  storesToCheck_2_15; // @[LoadQueue.scala 131:10:@9190.4]
  wire  storesToCheck_3_0; // @[LoadQueue.scala 131:10:@9232.4]
  wire  _T_8392; // @[LoadQueue.scala 131:81:@9235.4]
  wire  _T_8393; // @[LoadQueue.scala 131:72:@9236.4]
  wire  _T_8395; // @[LoadQueue.scala 132:33:@9237.4]
  wire  _T_8398; // @[LoadQueue.scala 132:41:@9239.4]
  wire  _T_8400; // @[LoadQueue.scala 132:9:@9240.4]
  wire  storesToCheck_3_1; // @[LoadQueue.scala 131:10:@9241.4]
  wire  _T_8406; // @[LoadQueue.scala 131:81:@9244.4]
  wire  _T_8407; // @[LoadQueue.scala 131:72:@9245.4]
  wire  _T_8409; // @[LoadQueue.scala 132:33:@9246.4]
  wire  _T_8412; // @[LoadQueue.scala 132:41:@9248.4]
  wire  _T_8414; // @[LoadQueue.scala 132:9:@9249.4]
  wire  storesToCheck_3_2; // @[LoadQueue.scala 131:10:@9250.4]
  wire  _T_8420; // @[LoadQueue.scala 131:81:@9253.4]
  wire  _T_8421; // @[LoadQueue.scala 131:72:@9254.4]
  wire  _T_8423; // @[LoadQueue.scala 132:33:@9255.4]
  wire  _T_8426; // @[LoadQueue.scala 132:41:@9257.4]
  wire  _T_8428; // @[LoadQueue.scala 132:9:@9258.4]
  wire  storesToCheck_3_3; // @[LoadQueue.scala 131:10:@9259.4]
  wire  _T_8434; // @[LoadQueue.scala 131:81:@9262.4]
  wire  _T_8435; // @[LoadQueue.scala 131:72:@9263.4]
  wire  _T_8437; // @[LoadQueue.scala 132:33:@9264.4]
  wire  _T_8440; // @[LoadQueue.scala 132:41:@9266.4]
  wire  _T_8442; // @[LoadQueue.scala 132:9:@9267.4]
  wire  storesToCheck_3_4; // @[LoadQueue.scala 131:10:@9268.4]
  wire  _T_8448; // @[LoadQueue.scala 131:81:@9271.4]
  wire  _T_8449; // @[LoadQueue.scala 131:72:@9272.4]
  wire  _T_8451; // @[LoadQueue.scala 132:33:@9273.4]
  wire  _T_8454; // @[LoadQueue.scala 132:41:@9275.4]
  wire  _T_8456; // @[LoadQueue.scala 132:9:@9276.4]
  wire  storesToCheck_3_5; // @[LoadQueue.scala 131:10:@9277.4]
  wire  _T_8462; // @[LoadQueue.scala 131:81:@9280.4]
  wire  _T_8463; // @[LoadQueue.scala 131:72:@9281.4]
  wire  _T_8465; // @[LoadQueue.scala 132:33:@9282.4]
  wire  _T_8468; // @[LoadQueue.scala 132:41:@9284.4]
  wire  _T_8470; // @[LoadQueue.scala 132:9:@9285.4]
  wire  storesToCheck_3_6; // @[LoadQueue.scala 131:10:@9286.4]
  wire  _T_8476; // @[LoadQueue.scala 131:81:@9289.4]
  wire  _T_8477; // @[LoadQueue.scala 131:72:@9290.4]
  wire  _T_8479; // @[LoadQueue.scala 132:33:@9291.4]
  wire  _T_8482; // @[LoadQueue.scala 132:41:@9293.4]
  wire  _T_8484; // @[LoadQueue.scala 132:9:@9294.4]
  wire  storesToCheck_3_7; // @[LoadQueue.scala 131:10:@9295.4]
  wire  _T_8490; // @[LoadQueue.scala 131:81:@9298.4]
  wire  _T_8491; // @[LoadQueue.scala 131:72:@9299.4]
  wire  _T_8493; // @[LoadQueue.scala 132:33:@9300.4]
  wire  _T_8496; // @[LoadQueue.scala 132:41:@9302.4]
  wire  _T_8498; // @[LoadQueue.scala 132:9:@9303.4]
  wire  storesToCheck_3_8; // @[LoadQueue.scala 131:10:@9304.4]
  wire  _T_8504; // @[LoadQueue.scala 131:81:@9307.4]
  wire  _T_8505; // @[LoadQueue.scala 131:72:@9308.4]
  wire  _T_8507; // @[LoadQueue.scala 132:33:@9309.4]
  wire  _T_8510; // @[LoadQueue.scala 132:41:@9311.4]
  wire  _T_8512; // @[LoadQueue.scala 132:9:@9312.4]
  wire  storesToCheck_3_9; // @[LoadQueue.scala 131:10:@9313.4]
  wire  _T_8518; // @[LoadQueue.scala 131:81:@9316.4]
  wire  _T_8519; // @[LoadQueue.scala 131:72:@9317.4]
  wire  _T_8521; // @[LoadQueue.scala 132:33:@9318.4]
  wire  _T_8524; // @[LoadQueue.scala 132:41:@9320.4]
  wire  _T_8526; // @[LoadQueue.scala 132:9:@9321.4]
  wire  storesToCheck_3_10; // @[LoadQueue.scala 131:10:@9322.4]
  wire  _T_8532; // @[LoadQueue.scala 131:81:@9325.4]
  wire  _T_8533; // @[LoadQueue.scala 131:72:@9326.4]
  wire  _T_8535; // @[LoadQueue.scala 132:33:@9327.4]
  wire  _T_8538; // @[LoadQueue.scala 132:41:@9329.4]
  wire  _T_8540; // @[LoadQueue.scala 132:9:@9330.4]
  wire  storesToCheck_3_11; // @[LoadQueue.scala 131:10:@9331.4]
  wire  _T_8546; // @[LoadQueue.scala 131:81:@9334.4]
  wire  _T_8547; // @[LoadQueue.scala 131:72:@9335.4]
  wire  _T_8549; // @[LoadQueue.scala 132:33:@9336.4]
  wire  _T_8552; // @[LoadQueue.scala 132:41:@9338.4]
  wire  _T_8554; // @[LoadQueue.scala 132:9:@9339.4]
  wire  storesToCheck_3_12; // @[LoadQueue.scala 131:10:@9340.4]
  wire  _T_8560; // @[LoadQueue.scala 131:81:@9343.4]
  wire  _T_8561; // @[LoadQueue.scala 131:72:@9344.4]
  wire  _T_8563; // @[LoadQueue.scala 132:33:@9345.4]
  wire  _T_8566; // @[LoadQueue.scala 132:41:@9347.4]
  wire  _T_8568; // @[LoadQueue.scala 132:9:@9348.4]
  wire  storesToCheck_3_13; // @[LoadQueue.scala 131:10:@9349.4]
  wire  _T_8574; // @[LoadQueue.scala 131:81:@9352.4]
  wire  _T_8575; // @[LoadQueue.scala 131:72:@9353.4]
  wire  _T_8577; // @[LoadQueue.scala 132:33:@9354.4]
  wire  _T_8580; // @[LoadQueue.scala 132:41:@9356.4]
  wire  _T_8582; // @[LoadQueue.scala 132:9:@9357.4]
  wire  storesToCheck_3_14; // @[LoadQueue.scala 131:10:@9358.4]
  wire  _T_8588; // @[LoadQueue.scala 131:81:@9361.4]
  wire  storesToCheck_3_15; // @[LoadQueue.scala 131:10:@9367.4]
  wire  storesToCheck_4_0; // @[LoadQueue.scala 131:10:@9409.4]
  wire  _T_8638; // @[LoadQueue.scala 131:81:@9412.4]
  wire  _T_8639; // @[LoadQueue.scala 131:72:@9413.4]
  wire  _T_8641; // @[LoadQueue.scala 132:33:@9414.4]
  wire  _T_8644; // @[LoadQueue.scala 132:41:@9416.4]
  wire  _T_8646; // @[LoadQueue.scala 132:9:@9417.4]
  wire  storesToCheck_4_1; // @[LoadQueue.scala 131:10:@9418.4]
  wire  _T_8652; // @[LoadQueue.scala 131:81:@9421.4]
  wire  _T_8653; // @[LoadQueue.scala 131:72:@9422.4]
  wire  _T_8655; // @[LoadQueue.scala 132:33:@9423.4]
  wire  _T_8658; // @[LoadQueue.scala 132:41:@9425.4]
  wire  _T_8660; // @[LoadQueue.scala 132:9:@9426.4]
  wire  storesToCheck_4_2; // @[LoadQueue.scala 131:10:@9427.4]
  wire  _T_8666; // @[LoadQueue.scala 131:81:@9430.4]
  wire  _T_8667; // @[LoadQueue.scala 131:72:@9431.4]
  wire  _T_8669; // @[LoadQueue.scala 132:33:@9432.4]
  wire  _T_8672; // @[LoadQueue.scala 132:41:@9434.4]
  wire  _T_8674; // @[LoadQueue.scala 132:9:@9435.4]
  wire  storesToCheck_4_3; // @[LoadQueue.scala 131:10:@9436.4]
  wire  _T_8680; // @[LoadQueue.scala 131:81:@9439.4]
  wire  _T_8681; // @[LoadQueue.scala 131:72:@9440.4]
  wire  _T_8683; // @[LoadQueue.scala 132:33:@9441.4]
  wire  _T_8686; // @[LoadQueue.scala 132:41:@9443.4]
  wire  _T_8688; // @[LoadQueue.scala 132:9:@9444.4]
  wire  storesToCheck_4_4; // @[LoadQueue.scala 131:10:@9445.4]
  wire  _T_8694; // @[LoadQueue.scala 131:81:@9448.4]
  wire  _T_8695; // @[LoadQueue.scala 131:72:@9449.4]
  wire  _T_8697; // @[LoadQueue.scala 132:33:@9450.4]
  wire  _T_8700; // @[LoadQueue.scala 132:41:@9452.4]
  wire  _T_8702; // @[LoadQueue.scala 132:9:@9453.4]
  wire  storesToCheck_4_5; // @[LoadQueue.scala 131:10:@9454.4]
  wire  _T_8708; // @[LoadQueue.scala 131:81:@9457.4]
  wire  _T_8709; // @[LoadQueue.scala 131:72:@9458.4]
  wire  _T_8711; // @[LoadQueue.scala 132:33:@9459.4]
  wire  _T_8714; // @[LoadQueue.scala 132:41:@9461.4]
  wire  _T_8716; // @[LoadQueue.scala 132:9:@9462.4]
  wire  storesToCheck_4_6; // @[LoadQueue.scala 131:10:@9463.4]
  wire  _T_8722; // @[LoadQueue.scala 131:81:@9466.4]
  wire  _T_8723; // @[LoadQueue.scala 131:72:@9467.4]
  wire  _T_8725; // @[LoadQueue.scala 132:33:@9468.4]
  wire  _T_8728; // @[LoadQueue.scala 132:41:@9470.4]
  wire  _T_8730; // @[LoadQueue.scala 132:9:@9471.4]
  wire  storesToCheck_4_7; // @[LoadQueue.scala 131:10:@9472.4]
  wire  _T_8736; // @[LoadQueue.scala 131:81:@9475.4]
  wire  _T_8737; // @[LoadQueue.scala 131:72:@9476.4]
  wire  _T_8739; // @[LoadQueue.scala 132:33:@9477.4]
  wire  _T_8742; // @[LoadQueue.scala 132:41:@9479.4]
  wire  _T_8744; // @[LoadQueue.scala 132:9:@9480.4]
  wire  storesToCheck_4_8; // @[LoadQueue.scala 131:10:@9481.4]
  wire  _T_8750; // @[LoadQueue.scala 131:81:@9484.4]
  wire  _T_8751; // @[LoadQueue.scala 131:72:@9485.4]
  wire  _T_8753; // @[LoadQueue.scala 132:33:@9486.4]
  wire  _T_8756; // @[LoadQueue.scala 132:41:@9488.4]
  wire  _T_8758; // @[LoadQueue.scala 132:9:@9489.4]
  wire  storesToCheck_4_9; // @[LoadQueue.scala 131:10:@9490.4]
  wire  _T_8764; // @[LoadQueue.scala 131:81:@9493.4]
  wire  _T_8765; // @[LoadQueue.scala 131:72:@9494.4]
  wire  _T_8767; // @[LoadQueue.scala 132:33:@9495.4]
  wire  _T_8770; // @[LoadQueue.scala 132:41:@9497.4]
  wire  _T_8772; // @[LoadQueue.scala 132:9:@9498.4]
  wire  storesToCheck_4_10; // @[LoadQueue.scala 131:10:@9499.4]
  wire  _T_8778; // @[LoadQueue.scala 131:81:@9502.4]
  wire  _T_8779; // @[LoadQueue.scala 131:72:@9503.4]
  wire  _T_8781; // @[LoadQueue.scala 132:33:@9504.4]
  wire  _T_8784; // @[LoadQueue.scala 132:41:@9506.4]
  wire  _T_8786; // @[LoadQueue.scala 132:9:@9507.4]
  wire  storesToCheck_4_11; // @[LoadQueue.scala 131:10:@9508.4]
  wire  _T_8792; // @[LoadQueue.scala 131:81:@9511.4]
  wire  _T_8793; // @[LoadQueue.scala 131:72:@9512.4]
  wire  _T_8795; // @[LoadQueue.scala 132:33:@9513.4]
  wire  _T_8798; // @[LoadQueue.scala 132:41:@9515.4]
  wire  _T_8800; // @[LoadQueue.scala 132:9:@9516.4]
  wire  storesToCheck_4_12; // @[LoadQueue.scala 131:10:@9517.4]
  wire  _T_8806; // @[LoadQueue.scala 131:81:@9520.4]
  wire  _T_8807; // @[LoadQueue.scala 131:72:@9521.4]
  wire  _T_8809; // @[LoadQueue.scala 132:33:@9522.4]
  wire  _T_8812; // @[LoadQueue.scala 132:41:@9524.4]
  wire  _T_8814; // @[LoadQueue.scala 132:9:@9525.4]
  wire  storesToCheck_4_13; // @[LoadQueue.scala 131:10:@9526.4]
  wire  _T_8820; // @[LoadQueue.scala 131:81:@9529.4]
  wire  _T_8821; // @[LoadQueue.scala 131:72:@9530.4]
  wire  _T_8823; // @[LoadQueue.scala 132:33:@9531.4]
  wire  _T_8826; // @[LoadQueue.scala 132:41:@9533.4]
  wire  _T_8828; // @[LoadQueue.scala 132:9:@9534.4]
  wire  storesToCheck_4_14; // @[LoadQueue.scala 131:10:@9535.4]
  wire  _T_8834; // @[LoadQueue.scala 131:81:@9538.4]
  wire  storesToCheck_4_15; // @[LoadQueue.scala 131:10:@9544.4]
  wire  storesToCheck_5_0; // @[LoadQueue.scala 131:10:@9586.4]
  wire  _T_8884; // @[LoadQueue.scala 131:81:@9589.4]
  wire  _T_8885; // @[LoadQueue.scala 131:72:@9590.4]
  wire  _T_8887; // @[LoadQueue.scala 132:33:@9591.4]
  wire  _T_8890; // @[LoadQueue.scala 132:41:@9593.4]
  wire  _T_8892; // @[LoadQueue.scala 132:9:@9594.4]
  wire  storesToCheck_5_1; // @[LoadQueue.scala 131:10:@9595.4]
  wire  _T_8898; // @[LoadQueue.scala 131:81:@9598.4]
  wire  _T_8899; // @[LoadQueue.scala 131:72:@9599.4]
  wire  _T_8901; // @[LoadQueue.scala 132:33:@9600.4]
  wire  _T_8904; // @[LoadQueue.scala 132:41:@9602.4]
  wire  _T_8906; // @[LoadQueue.scala 132:9:@9603.4]
  wire  storesToCheck_5_2; // @[LoadQueue.scala 131:10:@9604.4]
  wire  _T_8912; // @[LoadQueue.scala 131:81:@9607.4]
  wire  _T_8913; // @[LoadQueue.scala 131:72:@9608.4]
  wire  _T_8915; // @[LoadQueue.scala 132:33:@9609.4]
  wire  _T_8918; // @[LoadQueue.scala 132:41:@9611.4]
  wire  _T_8920; // @[LoadQueue.scala 132:9:@9612.4]
  wire  storesToCheck_5_3; // @[LoadQueue.scala 131:10:@9613.4]
  wire  _T_8926; // @[LoadQueue.scala 131:81:@9616.4]
  wire  _T_8927; // @[LoadQueue.scala 131:72:@9617.4]
  wire  _T_8929; // @[LoadQueue.scala 132:33:@9618.4]
  wire  _T_8932; // @[LoadQueue.scala 132:41:@9620.4]
  wire  _T_8934; // @[LoadQueue.scala 132:9:@9621.4]
  wire  storesToCheck_5_4; // @[LoadQueue.scala 131:10:@9622.4]
  wire  _T_8940; // @[LoadQueue.scala 131:81:@9625.4]
  wire  _T_8941; // @[LoadQueue.scala 131:72:@9626.4]
  wire  _T_8943; // @[LoadQueue.scala 132:33:@9627.4]
  wire  _T_8946; // @[LoadQueue.scala 132:41:@9629.4]
  wire  _T_8948; // @[LoadQueue.scala 132:9:@9630.4]
  wire  storesToCheck_5_5; // @[LoadQueue.scala 131:10:@9631.4]
  wire  _T_8954; // @[LoadQueue.scala 131:81:@9634.4]
  wire  _T_8955; // @[LoadQueue.scala 131:72:@9635.4]
  wire  _T_8957; // @[LoadQueue.scala 132:33:@9636.4]
  wire  _T_8960; // @[LoadQueue.scala 132:41:@9638.4]
  wire  _T_8962; // @[LoadQueue.scala 132:9:@9639.4]
  wire  storesToCheck_5_6; // @[LoadQueue.scala 131:10:@9640.4]
  wire  _T_8968; // @[LoadQueue.scala 131:81:@9643.4]
  wire  _T_8969; // @[LoadQueue.scala 131:72:@9644.4]
  wire  _T_8971; // @[LoadQueue.scala 132:33:@9645.4]
  wire  _T_8974; // @[LoadQueue.scala 132:41:@9647.4]
  wire  _T_8976; // @[LoadQueue.scala 132:9:@9648.4]
  wire  storesToCheck_5_7; // @[LoadQueue.scala 131:10:@9649.4]
  wire  _T_8982; // @[LoadQueue.scala 131:81:@9652.4]
  wire  _T_8983; // @[LoadQueue.scala 131:72:@9653.4]
  wire  _T_8985; // @[LoadQueue.scala 132:33:@9654.4]
  wire  _T_8988; // @[LoadQueue.scala 132:41:@9656.4]
  wire  _T_8990; // @[LoadQueue.scala 132:9:@9657.4]
  wire  storesToCheck_5_8; // @[LoadQueue.scala 131:10:@9658.4]
  wire  _T_8996; // @[LoadQueue.scala 131:81:@9661.4]
  wire  _T_8997; // @[LoadQueue.scala 131:72:@9662.4]
  wire  _T_8999; // @[LoadQueue.scala 132:33:@9663.4]
  wire  _T_9002; // @[LoadQueue.scala 132:41:@9665.4]
  wire  _T_9004; // @[LoadQueue.scala 132:9:@9666.4]
  wire  storesToCheck_5_9; // @[LoadQueue.scala 131:10:@9667.4]
  wire  _T_9010; // @[LoadQueue.scala 131:81:@9670.4]
  wire  _T_9011; // @[LoadQueue.scala 131:72:@9671.4]
  wire  _T_9013; // @[LoadQueue.scala 132:33:@9672.4]
  wire  _T_9016; // @[LoadQueue.scala 132:41:@9674.4]
  wire  _T_9018; // @[LoadQueue.scala 132:9:@9675.4]
  wire  storesToCheck_5_10; // @[LoadQueue.scala 131:10:@9676.4]
  wire  _T_9024; // @[LoadQueue.scala 131:81:@9679.4]
  wire  _T_9025; // @[LoadQueue.scala 131:72:@9680.4]
  wire  _T_9027; // @[LoadQueue.scala 132:33:@9681.4]
  wire  _T_9030; // @[LoadQueue.scala 132:41:@9683.4]
  wire  _T_9032; // @[LoadQueue.scala 132:9:@9684.4]
  wire  storesToCheck_5_11; // @[LoadQueue.scala 131:10:@9685.4]
  wire  _T_9038; // @[LoadQueue.scala 131:81:@9688.4]
  wire  _T_9039; // @[LoadQueue.scala 131:72:@9689.4]
  wire  _T_9041; // @[LoadQueue.scala 132:33:@9690.4]
  wire  _T_9044; // @[LoadQueue.scala 132:41:@9692.4]
  wire  _T_9046; // @[LoadQueue.scala 132:9:@9693.4]
  wire  storesToCheck_5_12; // @[LoadQueue.scala 131:10:@9694.4]
  wire  _T_9052; // @[LoadQueue.scala 131:81:@9697.4]
  wire  _T_9053; // @[LoadQueue.scala 131:72:@9698.4]
  wire  _T_9055; // @[LoadQueue.scala 132:33:@9699.4]
  wire  _T_9058; // @[LoadQueue.scala 132:41:@9701.4]
  wire  _T_9060; // @[LoadQueue.scala 132:9:@9702.4]
  wire  storesToCheck_5_13; // @[LoadQueue.scala 131:10:@9703.4]
  wire  _T_9066; // @[LoadQueue.scala 131:81:@9706.4]
  wire  _T_9067; // @[LoadQueue.scala 131:72:@9707.4]
  wire  _T_9069; // @[LoadQueue.scala 132:33:@9708.4]
  wire  _T_9072; // @[LoadQueue.scala 132:41:@9710.4]
  wire  _T_9074; // @[LoadQueue.scala 132:9:@9711.4]
  wire  storesToCheck_5_14; // @[LoadQueue.scala 131:10:@9712.4]
  wire  _T_9080; // @[LoadQueue.scala 131:81:@9715.4]
  wire  storesToCheck_5_15; // @[LoadQueue.scala 131:10:@9721.4]
  wire  storesToCheck_6_0; // @[LoadQueue.scala 131:10:@9763.4]
  wire  _T_9130; // @[LoadQueue.scala 131:81:@9766.4]
  wire  _T_9131; // @[LoadQueue.scala 131:72:@9767.4]
  wire  _T_9133; // @[LoadQueue.scala 132:33:@9768.4]
  wire  _T_9136; // @[LoadQueue.scala 132:41:@9770.4]
  wire  _T_9138; // @[LoadQueue.scala 132:9:@9771.4]
  wire  storesToCheck_6_1; // @[LoadQueue.scala 131:10:@9772.4]
  wire  _T_9144; // @[LoadQueue.scala 131:81:@9775.4]
  wire  _T_9145; // @[LoadQueue.scala 131:72:@9776.4]
  wire  _T_9147; // @[LoadQueue.scala 132:33:@9777.4]
  wire  _T_9150; // @[LoadQueue.scala 132:41:@9779.4]
  wire  _T_9152; // @[LoadQueue.scala 132:9:@9780.4]
  wire  storesToCheck_6_2; // @[LoadQueue.scala 131:10:@9781.4]
  wire  _T_9158; // @[LoadQueue.scala 131:81:@9784.4]
  wire  _T_9159; // @[LoadQueue.scala 131:72:@9785.4]
  wire  _T_9161; // @[LoadQueue.scala 132:33:@9786.4]
  wire  _T_9164; // @[LoadQueue.scala 132:41:@9788.4]
  wire  _T_9166; // @[LoadQueue.scala 132:9:@9789.4]
  wire  storesToCheck_6_3; // @[LoadQueue.scala 131:10:@9790.4]
  wire  _T_9172; // @[LoadQueue.scala 131:81:@9793.4]
  wire  _T_9173; // @[LoadQueue.scala 131:72:@9794.4]
  wire  _T_9175; // @[LoadQueue.scala 132:33:@9795.4]
  wire  _T_9178; // @[LoadQueue.scala 132:41:@9797.4]
  wire  _T_9180; // @[LoadQueue.scala 132:9:@9798.4]
  wire  storesToCheck_6_4; // @[LoadQueue.scala 131:10:@9799.4]
  wire  _T_9186; // @[LoadQueue.scala 131:81:@9802.4]
  wire  _T_9187; // @[LoadQueue.scala 131:72:@9803.4]
  wire  _T_9189; // @[LoadQueue.scala 132:33:@9804.4]
  wire  _T_9192; // @[LoadQueue.scala 132:41:@9806.4]
  wire  _T_9194; // @[LoadQueue.scala 132:9:@9807.4]
  wire  storesToCheck_6_5; // @[LoadQueue.scala 131:10:@9808.4]
  wire  _T_9200; // @[LoadQueue.scala 131:81:@9811.4]
  wire  _T_9201; // @[LoadQueue.scala 131:72:@9812.4]
  wire  _T_9203; // @[LoadQueue.scala 132:33:@9813.4]
  wire  _T_9206; // @[LoadQueue.scala 132:41:@9815.4]
  wire  _T_9208; // @[LoadQueue.scala 132:9:@9816.4]
  wire  storesToCheck_6_6; // @[LoadQueue.scala 131:10:@9817.4]
  wire  _T_9214; // @[LoadQueue.scala 131:81:@9820.4]
  wire  _T_9215; // @[LoadQueue.scala 131:72:@9821.4]
  wire  _T_9217; // @[LoadQueue.scala 132:33:@9822.4]
  wire  _T_9220; // @[LoadQueue.scala 132:41:@9824.4]
  wire  _T_9222; // @[LoadQueue.scala 132:9:@9825.4]
  wire  storesToCheck_6_7; // @[LoadQueue.scala 131:10:@9826.4]
  wire  _T_9228; // @[LoadQueue.scala 131:81:@9829.4]
  wire  _T_9229; // @[LoadQueue.scala 131:72:@9830.4]
  wire  _T_9231; // @[LoadQueue.scala 132:33:@9831.4]
  wire  _T_9234; // @[LoadQueue.scala 132:41:@9833.4]
  wire  _T_9236; // @[LoadQueue.scala 132:9:@9834.4]
  wire  storesToCheck_6_8; // @[LoadQueue.scala 131:10:@9835.4]
  wire  _T_9242; // @[LoadQueue.scala 131:81:@9838.4]
  wire  _T_9243; // @[LoadQueue.scala 131:72:@9839.4]
  wire  _T_9245; // @[LoadQueue.scala 132:33:@9840.4]
  wire  _T_9248; // @[LoadQueue.scala 132:41:@9842.4]
  wire  _T_9250; // @[LoadQueue.scala 132:9:@9843.4]
  wire  storesToCheck_6_9; // @[LoadQueue.scala 131:10:@9844.4]
  wire  _T_9256; // @[LoadQueue.scala 131:81:@9847.4]
  wire  _T_9257; // @[LoadQueue.scala 131:72:@9848.4]
  wire  _T_9259; // @[LoadQueue.scala 132:33:@9849.4]
  wire  _T_9262; // @[LoadQueue.scala 132:41:@9851.4]
  wire  _T_9264; // @[LoadQueue.scala 132:9:@9852.4]
  wire  storesToCheck_6_10; // @[LoadQueue.scala 131:10:@9853.4]
  wire  _T_9270; // @[LoadQueue.scala 131:81:@9856.4]
  wire  _T_9271; // @[LoadQueue.scala 131:72:@9857.4]
  wire  _T_9273; // @[LoadQueue.scala 132:33:@9858.4]
  wire  _T_9276; // @[LoadQueue.scala 132:41:@9860.4]
  wire  _T_9278; // @[LoadQueue.scala 132:9:@9861.4]
  wire  storesToCheck_6_11; // @[LoadQueue.scala 131:10:@9862.4]
  wire  _T_9284; // @[LoadQueue.scala 131:81:@9865.4]
  wire  _T_9285; // @[LoadQueue.scala 131:72:@9866.4]
  wire  _T_9287; // @[LoadQueue.scala 132:33:@9867.4]
  wire  _T_9290; // @[LoadQueue.scala 132:41:@9869.4]
  wire  _T_9292; // @[LoadQueue.scala 132:9:@9870.4]
  wire  storesToCheck_6_12; // @[LoadQueue.scala 131:10:@9871.4]
  wire  _T_9298; // @[LoadQueue.scala 131:81:@9874.4]
  wire  _T_9299; // @[LoadQueue.scala 131:72:@9875.4]
  wire  _T_9301; // @[LoadQueue.scala 132:33:@9876.4]
  wire  _T_9304; // @[LoadQueue.scala 132:41:@9878.4]
  wire  _T_9306; // @[LoadQueue.scala 132:9:@9879.4]
  wire  storesToCheck_6_13; // @[LoadQueue.scala 131:10:@9880.4]
  wire  _T_9312; // @[LoadQueue.scala 131:81:@9883.4]
  wire  _T_9313; // @[LoadQueue.scala 131:72:@9884.4]
  wire  _T_9315; // @[LoadQueue.scala 132:33:@9885.4]
  wire  _T_9318; // @[LoadQueue.scala 132:41:@9887.4]
  wire  _T_9320; // @[LoadQueue.scala 132:9:@9888.4]
  wire  storesToCheck_6_14; // @[LoadQueue.scala 131:10:@9889.4]
  wire  _T_9326; // @[LoadQueue.scala 131:81:@9892.4]
  wire  storesToCheck_6_15; // @[LoadQueue.scala 131:10:@9898.4]
  wire  storesToCheck_7_0; // @[LoadQueue.scala 131:10:@9940.4]
  wire  _T_9376; // @[LoadQueue.scala 131:81:@9943.4]
  wire  _T_9377; // @[LoadQueue.scala 131:72:@9944.4]
  wire  _T_9379; // @[LoadQueue.scala 132:33:@9945.4]
  wire  _T_9382; // @[LoadQueue.scala 132:41:@9947.4]
  wire  _T_9384; // @[LoadQueue.scala 132:9:@9948.4]
  wire  storesToCheck_7_1; // @[LoadQueue.scala 131:10:@9949.4]
  wire  _T_9390; // @[LoadQueue.scala 131:81:@9952.4]
  wire  _T_9391; // @[LoadQueue.scala 131:72:@9953.4]
  wire  _T_9393; // @[LoadQueue.scala 132:33:@9954.4]
  wire  _T_9396; // @[LoadQueue.scala 132:41:@9956.4]
  wire  _T_9398; // @[LoadQueue.scala 132:9:@9957.4]
  wire  storesToCheck_7_2; // @[LoadQueue.scala 131:10:@9958.4]
  wire  _T_9404; // @[LoadQueue.scala 131:81:@9961.4]
  wire  _T_9405; // @[LoadQueue.scala 131:72:@9962.4]
  wire  _T_9407; // @[LoadQueue.scala 132:33:@9963.4]
  wire  _T_9410; // @[LoadQueue.scala 132:41:@9965.4]
  wire  _T_9412; // @[LoadQueue.scala 132:9:@9966.4]
  wire  storesToCheck_7_3; // @[LoadQueue.scala 131:10:@9967.4]
  wire  _T_9418; // @[LoadQueue.scala 131:81:@9970.4]
  wire  _T_9419; // @[LoadQueue.scala 131:72:@9971.4]
  wire  _T_9421; // @[LoadQueue.scala 132:33:@9972.4]
  wire  _T_9424; // @[LoadQueue.scala 132:41:@9974.4]
  wire  _T_9426; // @[LoadQueue.scala 132:9:@9975.4]
  wire  storesToCheck_7_4; // @[LoadQueue.scala 131:10:@9976.4]
  wire  _T_9432; // @[LoadQueue.scala 131:81:@9979.4]
  wire  _T_9433; // @[LoadQueue.scala 131:72:@9980.4]
  wire  _T_9435; // @[LoadQueue.scala 132:33:@9981.4]
  wire  _T_9438; // @[LoadQueue.scala 132:41:@9983.4]
  wire  _T_9440; // @[LoadQueue.scala 132:9:@9984.4]
  wire  storesToCheck_7_5; // @[LoadQueue.scala 131:10:@9985.4]
  wire  _T_9446; // @[LoadQueue.scala 131:81:@9988.4]
  wire  _T_9447; // @[LoadQueue.scala 131:72:@9989.4]
  wire  _T_9449; // @[LoadQueue.scala 132:33:@9990.4]
  wire  _T_9452; // @[LoadQueue.scala 132:41:@9992.4]
  wire  _T_9454; // @[LoadQueue.scala 132:9:@9993.4]
  wire  storesToCheck_7_6; // @[LoadQueue.scala 131:10:@9994.4]
  wire  _T_9460; // @[LoadQueue.scala 131:81:@9997.4]
  wire  _T_9461; // @[LoadQueue.scala 131:72:@9998.4]
  wire  _T_9463; // @[LoadQueue.scala 132:33:@9999.4]
  wire  _T_9466; // @[LoadQueue.scala 132:41:@10001.4]
  wire  _T_9468; // @[LoadQueue.scala 132:9:@10002.4]
  wire  storesToCheck_7_7; // @[LoadQueue.scala 131:10:@10003.4]
  wire  _T_9474; // @[LoadQueue.scala 131:81:@10006.4]
  wire  _T_9475; // @[LoadQueue.scala 131:72:@10007.4]
  wire  _T_9477; // @[LoadQueue.scala 132:33:@10008.4]
  wire  _T_9480; // @[LoadQueue.scala 132:41:@10010.4]
  wire  _T_9482; // @[LoadQueue.scala 132:9:@10011.4]
  wire  storesToCheck_7_8; // @[LoadQueue.scala 131:10:@10012.4]
  wire  _T_9488; // @[LoadQueue.scala 131:81:@10015.4]
  wire  _T_9489; // @[LoadQueue.scala 131:72:@10016.4]
  wire  _T_9491; // @[LoadQueue.scala 132:33:@10017.4]
  wire  _T_9494; // @[LoadQueue.scala 132:41:@10019.4]
  wire  _T_9496; // @[LoadQueue.scala 132:9:@10020.4]
  wire  storesToCheck_7_9; // @[LoadQueue.scala 131:10:@10021.4]
  wire  _T_9502; // @[LoadQueue.scala 131:81:@10024.4]
  wire  _T_9503; // @[LoadQueue.scala 131:72:@10025.4]
  wire  _T_9505; // @[LoadQueue.scala 132:33:@10026.4]
  wire  _T_9508; // @[LoadQueue.scala 132:41:@10028.4]
  wire  _T_9510; // @[LoadQueue.scala 132:9:@10029.4]
  wire  storesToCheck_7_10; // @[LoadQueue.scala 131:10:@10030.4]
  wire  _T_9516; // @[LoadQueue.scala 131:81:@10033.4]
  wire  _T_9517; // @[LoadQueue.scala 131:72:@10034.4]
  wire  _T_9519; // @[LoadQueue.scala 132:33:@10035.4]
  wire  _T_9522; // @[LoadQueue.scala 132:41:@10037.4]
  wire  _T_9524; // @[LoadQueue.scala 132:9:@10038.4]
  wire  storesToCheck_7_11; // @[LoadQueue.scala 131:10:@10039.4]
  wire  _T_9530; // @[LoadQueue.scala 131:81:@10042.4]
  wire  _T_9531; // @[LoadQueue.scala 131:72:@10043.4]
  wire  _T_9533; // @[LoadQueue.scala 132:33:@10044.4]
  wire  _T_9536; // @[LoadQueue.scala 132:41:@10046.4]
  wire  _T_9538; // @[LoadQueue.scala 132:9:@10047.4]
  wire  storesToCheck_7_12; // @[LoadQueue.scala 131:10:@10048.4]
  wire  _T_9544; // @[LoadQueue.scala 131:81:@10051.4]
  wire  _T_9545; // @[LoadQueue.scala 131:72:@10052.4]
  wire  _T_9547; // @[LoadQueue.scala 132:33:@10053.4]
  wire  _T_9550; // @[LoadQueue.scala 132:41:@10055.4]
  wire  _T_9552; // @[LoadQueue.scala 132:9:@10056.4]
  wire  storesToCheck_7_13; // @[LoadQueue.scala 131:10:@10057.4]
  wire  _T_9558; // @[LoadQueue.scala 131:81:@10060.4]
  wire  _T_9559; // @[LoadQueue.scala 131:72:@10061.4]
  wire  _T_9561; // @[LoadQueue.scala 132:33:@10062.4]
  wire  _T_9564; // @[LoadQueue.scala 132:41:@10064.4]
  wire  _T_9566; // @[LoadQueue.scala 132:9:@10065.4]
  wire  storesToCheck_7_14; // @[LoadQueue.scala 131:10:@10066.4]
  wire  _T_9572; // @[LoadQueue.scala 131:81:@10069.4]
  wire  storesToCheck_7_15; // @[LoadQueue.scala 131:10:@10075.4]
  wire  storesToCheck_8_0; // @[LoadQueue.scala 131:10:@10117.4]
  wire  _T_9622; // @[LoadQueue.scala 131:81:@10120.4]
  wire  _T_9623; // @[LoadQueue.scala 131:72:@10121.4]
  wire  _T_9625; // @[LoadQueue.scala 132:33:@10122.4]
  wire  _T_9628; // @[LoadQueue.scala 132:41:@10124.4]
  wire  _T_9630; // @[LoadQueue.scala 132:9:@10125.4]
  wire  storesToCheck_8_1; // @[LoadQueue.scala 131:10:@10126.4]
  wire  _T_9636; // @[LoadQueue.scala 131:81:@10129.4]
  wire  _T_9637; // @[LoadQueue.scala 131:72:@10130.4]
  wire  _T_9639; // @[LoadQueue.scala 132:33:@10131.4]
  wire  _T_9642; // @[LoadQueue.scala 132:41:@10133.4]
  wire  _T_9644; // @[LoadQueue.scala 132:9:@10134.4]
  wire  storesToCheck_8_2; // @[LoadQueue.scala 131:10:@10135.4]
  wire  _T_9650; // @[LoadQueue.scala 131:81:@10138.4]
  wire  _T_9651; // @[LoadQueue.scala 131:72:@10139.4]
  wire  _T_9653; // @[LoadQueue.scala 132:33:@10140.4]
  wire  _T_9656; // @[LoadQueue.scala 132:41:@10142.4]
  wire  _T_9658; // @[LoadQueue.scala 132:9:@10143.4]
  wire  storesToCheck_8_3; // @[LoadQueue.scala 131:10:@10144.4]
  wire  _T_9664; // @[LoadQueue.scala 131:81:@10147.4]
  wire  _T_9665; // @[LoadQueue.scala 131:72:@10148.4]
  wire  _T_9667; // @[LoadQueue.scala 132:33:@10149.4]
  wire  _T_9670; // @[LoadQueue.scala 132:41:@10151.4]
  wire  _T_9672; // @[LoadQueue.scala 132:9:@10152.4]
  wire  storesToCheck_8_4; // @[LoadQueue.scala 131:10:@10153.4]
  wire  _T_9678; // @[LoadQueue.scala 131:81:@10156.4]
  wire  _T_9679; // @[LoadQueue.scala 131:72:@10157.4]
  wire  _T_9681; // @[LoadQueue.scala 132:33:@10158.4]
  wire  _T_9684; // @[LoadQueue.scala 132:41:@10160.4]
  wire  _T_9686; // @[LoadQueue.scala 132:9:@10161.4]
  wire  storesToCheck_8_5; // @[LoadQueue.scala 131:10:@10162.4]
  wire  _T_9692; // @[LoadQueue.scala 131:81:@10165.4]
  wire  _T_9693; // @[LoadQueue.scala 131:72:@10166.4]
  wire  _T_9695; // @[LoadQueue.scala 132:33:@10167.4]
  wire  _T_9698; // @[LoadQueue.scala 132:41:@10169.4]
  wire  _T_9700; // @[LoadQueue.scala 132:9:@10170.4]
  wire  storesToCheck_8_6; // @[LoadQueue.scala 131:10:@10171.4]
  wire  _T_9706; // @[LoadQueue.scala 131:81:@10174.4]
  wire  _T_9707; // @[LoadQueue.scala 131:72:@10175.4]
  wire  _T_9709; // @[LoadQueue.scala 132:33:@10176.4]
  wire  _T_9712; // @[LoadQueue.scala 132:41:@10178.4]
  wire  _T_9714; // @[LoadQueue.scala 132:9:@10179.4]
  wire  storesToCheck_8_7; // @[LoadQueue.scala 131:10:@10180.4]
  wire  _T_9720; // @[LoadQueue.scala 131:81:@10183.4]
  wire  _T_9721; // @[LoadQueue.scala 131:72:@10184.4]
  wire  _T_9723; // @[LoadQueue.scala 132:33:@10185.4]
  wire  _T_9726; // @[LoadQueue.scala 132:41:@10187.4]
  wire  _T_9728; // @[LoadQueue.scala 132:9:@10188.4]
  wire  storesToCheck_8_8; // @[LoadQueue.scala 131:10:@10189.4]
  wire  _T_9734; // @[LoadQueue.scala 131:81:@10192.4]
  wire  _T_9735; // @[LoadQueue.scala 131:72:@10193.4]
  wire  _T_9737; // @[LoadQueue.scala 132:33:@10194.4]
  wire  _T_9740; // @[LoadQueue.scala 132:41:@10196.4]
  wire  _T_9742; // @[LoadQueue.scala 132:9:@10197.4]
  wire  storesToCheck_8_9; // @[LoadQueue.scala 131:10:@10198.4]
  wire  _T_9748; // @[LoadQueue.scala 131:81:@10201.4]
  wire  _T_9749; // @[LoadQueue.scala 131:72:@10202.4]
  wire  _T_9751; // @[LoadQueue.scala 132:33:@10203.4]
  wire  _T_9754; // @[LoadQueue.scala 132:41:@10205.4]
  wire  _T_9756; // @[LoadQueue.scala 132:9:@10206.4]
  wire  storesToCheck_8_10; // @[LoadQueue.scala 131:10:@10207.4]
  wire  _T_9762; // @[LoadQueue.scala 131:81:@10210.4]
  wire  _T_9763; // @[LoadQueue.scala 131:72:@10211.4]
  wire  _T_9765; // @[LoadQueue.scala 132:33:@10212.4]
  wire  _T_9768; // @[LoadQueue.scala 132:41:@10214.4]
  wire  _T_9770; // @[LoadQueue.scala 132:9:@10215.4]
  wire  storesToCheck_8_11; // @[LoadQueue.scala 131:10:@10216.4]
  wire  _T_9776; // @[LoadQueue.scala 131:81:@10219.4]
  wire  _T_9777; // @[LoadQueue.scala 131:72:@10220.4]
  wire  _T_9779; // @[LoadQueue.scala 132:33:@10221.4]
  wire  _T_9782; // @[LoadQueue.scala 132:41:@10223.4]
  wire  _T_9784; // @[LoadQueue.scala 132:9:@10224.4]
  wire  storesToCheck_8_12; // @[LoadQueue.scala 131:10:@10225.4]
  wire  _T_9790; // @[LoadQueue.scala 131:81:@10228.4]
  wire  _T_9791; // @[LoadQueue.scala 131:72:@10229.4]
  wire  _T_9793; // @[LoadQueue.scala 132:33:@10230.4]
  wire  _T_9796; // @[LoadQueue.scala 132:41:@10232.4]
  wire  _T_9798; // @[LoadQueue.scala 132:9:@10233.4]
  wire  storesToCheck_8_13; // @[LoadQueue.scala 131:10:@10234.4]
  wire  _T_9804; // @[LoadQueue.scala 131:81:@10237.4]
  wire  _T_9805; // @[LoadQueue.scala 131:72:@10238.4]
  wire  _T_9807; // @[LoadQueue.scala 132:33:@10239.4]
  wire  _T_9810; // @[LoadQueue.scala 132:41:@10241.4]
  wire  _T_9812; // @[LoadQueue.scala 132:9:@10242.4]
  wire  storesToCheck_8_14; // @[LoadQueue.scala 131:10:@10243.4]
  wire  _T_9818; // @[LoadQueue.scala 131:81:@10246.4]
  wire  storesToCheck_8_15; // @[LoadQueue.scala 131:10:@10252.4]
  wire  storesToCheck_9_0; // @[LoadQueue.scala 131:10:@10294.4]
  wire  _T_9868; // @[LoadQueue.scala 131:81:@10297.4]
  wire  _T_9869; // @[LoadQueue.scala 131:72:@10298.4]
  wire  _T_9871; // @[LoadQueue.scala 132:33:@10299.4]
  wire  _T_9874; // @[LoadQueue.scala 132:41:@10301.4]
  wire  _T_9876; // @[LoadQueue.scala 132:9:@10302.4]
  wire  storesToCheck_9_1; // @[LoadQueue.scala 131:10:@10303.4]
  wire  _T_9882; // @[LoadQueue.scala 131:81:@10306.4]
  wire  _T_9883; // @[LoadQueue.scala 131:72:@10307.4]
  wire  _T_9885; // @[LoadQueue.scala 132:33:@10308.4]
  wire  _T_9888; // @[LoadQueue.scala 132:41:@10310.4]
  wire  _T_9890; // @[LoadQueue.scala 132:9:@10311.4]
  wire  storesToCheck_9_2; // @[LoadQueue.scala 131:10:@10312.4]
  wire  _T_9896; // @[LoadQueue.scala 131:81:@10315.4]
  wire  _T_9897; // @[LoadQueue.scala 131:72:@10316.4]
  wire  _T_9899; // @[LoadQueue.scala 132:33:@10317.4]
  wire  _T_9902; // @[LoadQueue.scala 132:41:@10319.4]
  wire  _T_9904; // @[LoadQueue.scala 132:9:@10320.4]
  wire  storesToCheck_9_3; // @[LoadQueue.scala 131:10:@10321.4]
  wire  _T_9910; // @[LoadQueue.scala 131:81:@10324.4]
  wire  _T_9911; // @[LoadQueue.scala 131:72:@10325.4]
  wire  _T_9913; // @[LoadQueue.scala 132:33:@10326.4]
  wire  _T_9916; // @[LoadQueue.scala 132:41:@10328.4]
  wire  _T_9918; // @[LoadQueue.scala 132:9:@10329.4]
  wire  storesToCheck_9_4; // @[LoadQueue.scala 131:10:@10330.4]
  wire  _T_9924; // @[LoadQueue.scala 131:81:@10333.4]
  wire  _T_9925; // @[LoadQueue.scala 131:72:@10334.4]
  wire  _T_9927; // @[LoadQueue.scala 132:33:@10335.4]
  wire  _T_9930; // @[LoadQueue.scala 132:41:@10337.4]
  wire  _T_9932; // @[LoadQueue.scala 132:9:@10338.4]
  wire  storesToCheck_9_5; // @[LoadQueue.scala 131:10:@10339.4]
  wire  _T_9938; // @[LoadQueue.scala 131:81:@10342.4]
  wire  _T_9939; // @[LoadQueue.scala 131:72:@10343.4]
  wire  _T_9941; // @[LoadQueue.scala 132:33:@10344.4]
  wire  _T_9944; // @[LoadQueue.scala 132:41:@10346.4]
  wire  _T_9946; // @[LoadQueue.scala 132:9:@10347.4]
  wire  storesToCheck_9_6; // @[LoadQueue.scala 131:10:@10348.4]
  wire  _T_9952; // @[LoadQueue.scala 131:81:@10351.4]
  wire  _T_9953; // @[LoadQueue.scala 131:72:@10352.4]
  wire  _T_9955; // @[LoadQueue.scala 132:33:@10353.4]
  wire  _T_9958; // @[LoadQueue.scala 132:41:@10355.4]
  wire  _T_9960; // @[LoadQueue.scala 132:9:@10356.4]
  wire  storesToCheck_9_7; // @[LoadQueue.scala 131:10:@10357.4]
  wire  _T_9966; // @[LoadQueue.scala 131:81:@10360.4]
  wire  _T_9967; // @[LoadQueue.scala 131:72:@10361.4]
  wire  _T_9969; // @[LoadQueue.scala 132:33:@10362.4]
  wire  _T_9972; // @[LoadQueue.scala 132:41:@10364.4]
  wire  _T_9974; // @[LoadQueue.scala 132:9:@10365.4]
  wire  storesToCheck_9_8; // @[LoadQueue.scala 131:10:@10366.4]
  wire  _T_9980; // @[LoadQueue.scala 131:81:@10369.4]
  wire  _T_9981; // @[LoadQueue.scala 131:72:@10370.4]
  wire  _T_9983; // @[LoadQueue.scala 132:33:@10371.4]
  wire  _T_9986; // @[LoadQueue.scala 132:41:@10373.4]
  wire  _T_9988; // @[LoadQueue.scala 132:9:@10374.4]
  wire  storesToCheck_9_9; // @[LoadQueue.scala 131:10:@10375.4]
  wire  _T_9994; // @[LoadQueue.scala 131:81:@10378.4]
  wire  _T_9995; // @[LoadQueue.scala 131:72:@10379.4]
  wire  _T_9997; // @[LoadQueue.scala 132:33:@10380.4]
  wire  _T_10000; // @[LoadQueue.scala 132:41:@10382.4]
  wire  _T_10002; // @[LoadQueue.scala 132:9:@10383.4]
  wire  storesToCheck_9_10; // @[LoadQueue.scala 131:10:@10384.4]
  wire  _T_10008; // @[LoadQueue.scala 131:81:@10387.4]
  wire  _T_10009; // @[LoadQueue.scala 131:72:@10388.4]
  wire  _T_10011; // @[LoadQueue.scala 132:33:@10389.4]
  wire  _T_10014; // @[LoadQueue.scala 132:41:@10391.4]
  wire  _T_10016; // @[LoadQueue.scala 132:9:@10392.4]
  wire  storesToCheck_9_11; // @[LoadQueue.scala 131:10:@10393.4]
  wire  _T_10022; // @[LoadQueue.scala 131:81:@10396.4]
  wire  _T_10023; // @[LoadQueue.scala 131:72:@10397.4]
  wire  _T_10025; // @[LoadQueue.scala 132:33:@10398.4]
  wire  _T_10028; // @[LoadQueue.scala 132:41:@10400.4]
  wire  _T_10030; // @[LoadQueue.scala 132:9:@10401.4]
  wire  storesToCheck_9_12; // @[LoadQueue.scala 131:10:@10402.4]
  wire  _T_10036; // @[LoadQueue.scala 131:81:@10405.4]
  wire  _T_10037; // @[LoadQueue.scala 131:72:@10406.4]
  wire  _T_10039; // @[LoadQueue.scala 132:33:@10407.4]
  wire  _T_10042; // @[LoadQueue.scala 132:41:@10409.4]
  wire  _T_10044; // @[LoadQueue.scala 132:9:@10410.4]
  wire  storesToCheck_9_13; // @[LoadQueue.scala 131:10:@10411.4]
  wire  _T_10050; // @[LoadQueue.scala 131:81:@10414.4]
  wire  _T_10051; // @[LoadQueue.scala 131:72:@10415.4]
  wire  _T_10053; // @[LoadQueue.scala 132:33:@10416.4]
  wire  _T_10056; // @[LoadQueue.scala 132:41:@10418.4]
  wire  _T_10058; // @[LoadQueue.scala 132:9:@10419.4]
  wire  storesToCheck_9_14; // @[LoadQueue.scala 131:10:@10420.4]
  wire  _T_10064; // @[LoadQueue.scala 131:81:@10423.4]
  wire  storesToCheck_9_15; // @[LoadQueue.scala 131:10:@10429.4]
  wire  storesToCheck_10_0; // @[LoadQueue.scala 131:10:@10471.4]
  wire  _T_10114; // @[LoadQueue.scala 131:81:@10474.4]
  wire  _T_10115; // @[LoadQueue.scala 131:72:@10475.4]
  wire  _T_10117; // @[LoadQueue.scala 132:33:@10476.4]
  wire  _T_10120; // @[LoadQueue.scala 132:41:@10478.4]
  wire  _T_10122; // @[LoadQueue.scala 132:9:@10479.4]
  wire  storesToCheck_10_1; // @[LoadQueue.scala 131:10:@10480.4]
  wire  _T_10128; // @[LoadQueue.scala 131:81:@10483.4]
  wire  _T_10129; // @[LoadQueue.scala 131:72:@10484.4]
  wire  _T_10131; // @[LoadQueue.scala 132:33:@10485.4]
  wire  _T_10134; // @[LoadQueue.scala 132:41:@10487.4]
  wire  _T_10136; // @[LoadQueue.scala 132:9:@10488.4]
  wire  storesToCheck_10_2; // @[LoadQueue.scala 131:10:@10489.4]
  wire  _T_10142; // @[LoadQueue.scala 131:81:@10492.4]
  wire  _T_10143; // @[LoadQueue.scala 131:72:@10493.4]
  wire  _T_10145; // @[LoadQueue.scala 132:33:@10494.4]
  wire  _T_10148; // @[LoadQueue.scala 132:41:@10496.4]
  wire  _T_10150; // @[LoadQueue.scala 132:9:@10497.4]
  wire  storesToCheck_10_3; // @[LoadQueue.scala 131:10:@10498.4]
  wire  _T_10156; // @[LoadQueue.scala 131:81:@10501.4]
  wire  _T_10157; // @[LoadQueue.scala 131:72:@10502.4]
  wire  _T_10159; // @[LoadQueue.scala 132:33:@10503.4]
  wire  _T_10162; // @[LoadQueue.scala 132:41:@10505.4]
  wire  _T_10164; // @[LoadQueue.scala 132:9:@10506.4]
  wire  storesToCheck_10_4; // @[LoadQueue.scala 131:10:@10507.4]
  wire  _T_10170; // @[LoadQueue.scala 131:81:@10510.4]
  wire  _T_10171; // @[LoadQueue.scala 131:72:@10511.4]
  wire  _T_10173; // @[LoadQueue.scala 132:33:@10512.4]
  wire  _T_10176; // @[LoadQueue.scala 132:41:@10514.4]
  wire  _T_10178; // @[LoadQueue.scala 132:9:@10515.4]
  wire  storesToCheck_10_5; // @[LoadQueue.scala 131:10:@10516.4]
  wire  _T_10184; // @[LoadQueue.scala 131:81:@10519.4]
  wire  _T_10185; // @[LoadQueue.scala 131:72:@10520.4]
  wire  _T_10187; // @[LoadQueue.scala 132:33:@10521.4]
  wire  _T_10190; // @[LoadQueue.scala 132:41:@10523.4]
  wire  _T_10192; // @[LoadQueue.scala 132:9:@10524.4]
  wire  storesToCheck_10_6; // @[LoadQueue.scala 131:10:@10525.4]
  wire  _T_10198; // @[LoadQueue.scala 131:81:@10528.4]
  wire  _T_10199; // @[LoadQueue.scala 131:72:@10529.4]
  wire  _T_10201; // @[LoadQueue.scala 132:33:@10530.4]
  wire  _T_10204; // @[LoadQueue.scala 132:41:@10532.4]
  wire  _T_10206; // @[LoadQueue.scala 132:9:@10533.4]
  wire  storesToCheck_10_7; // @[LoadQueue.scala 131:10:@10534.4]
  wire  _T_10212; // @[LoadQueue.scala 131:81:@10537.4]
  wire  _T_10213; // @[LoadQueue.scala 131:72:@10538.4]
  wire  _T_10215; // @[LoadQueue.scala 132:33:@10539.4]
  wire  _T_10218; // @[LoadQueue.scala 132:41:@10541.4]
  wire  _T_10220; // @[LoadQueue.scala 132:9:@10542.4]
  wire  storesToCheck_10_8; // @[LoadQueue.scala 131:10:@10543.4]
  wire  _T_10226; // @[LoadQueue.scala 131:81:@10546.4]
  wire  _T_10227; // @[LoadQueue.scala 131:72:@10547.4]
  wire  _T_10229; // @[LoadQueue.scala 132:33:@10548.4]
  wire  _T_10232; // @[LoadQueue.scala 132:41:@10550.4]
  wire  _T_10234; // @[LoadQueue.scala 132:9:@10551.4]
  wire  storesToCheck_10_9; // @[LoadQueue.scala 131:10:@10552.4]
  wire  _T_10240; // @[LoadQueue.scala 131:81:@10555.4]
  wire  _T_10241; // @[LoadQueue.scala 131:72:@10556.4]
  wire  _T_10243; // @[LoadQueue.scala 132:33:@10557.4]
  wire  _T_10246; // @[LoadQueue.scala 132:41:@10559.4]
  wire  _T_10248; // @[LoadQueue.scala 132:9:@10560.4]
  wire  storesToCheck_10_10; // @[LoadQueue.scala 131:10:@10561.4]
  wire  _T_10254; // @[LoadQueue.scala 131:81:@10564.4]
  wire  _T_10255; // @[LoadQueue.scala 131:72:@10565.4]
  wire  _T_10257; // @[LoadQueue.scala 132:33:@10566.4]
  wire  _T_10260; // @[LoadQueue.scala 132:41:@10568.4]
  wire  _T_10262; // @[LoadQueue.scala 132:9:@10569.4]
  wire  storesToCheck_10_11; // @[LoadQueue.scala 131:10:@10570.4]
  wire  _T_10268; // @[LoadQueue.scala 131:81:@10573.4]
  wire  _T_10269; // @[LoadQueue.scala 131:72:@10574.4]
  wire  _T_10271; // @[LoadQueue.scala 132:33:@10575.4]
  wire  _T_10274; // @[LoadQueue.scala 132:41:@10577.4]
  wire  _T_10276; // @[LoadQueue.scala 132:9:@10578.4]
  wire  storesToCheck_10_12; // @[LoadQueue.scala 131:10:@10579.4]
  wire  _T_10282; // @[LoadQueue.scala 131:81:@10582.4]
  wire  _T_10283; // @[LoadQueue.scala 131:72:@10583.4]
  wire  _T_10285; // @[LoadQueue.scala 132:33:@10584.4]
  wire  _T_10288; // @[LoadQueue.scala 132:41:@10586.4]
  wire  _T_10290; // @[LoadQueue.scala 132:9:@10587.4]
  wire  storesToCheck_10_13; // @[LoadQueue.scala 131:10:@10588.4]
  wire  _T_10296; // @[LoadQueue.scala 131:81:@10591.4]
  wire  _T_10297; // @[LoadQueue.scala 131:72:@10592.4]
  wire  _T_10299; // @[LoadQueue.scala 132:33:@10593.4]
  wire  _T_10302; // @[LoadQueue.scala 132:41:@10595.4]
  wire  _T_10304; // @[LoadQueue.scala 132:9:@10596.4]
  wire  storesToCheck_10_14; // @[LoadQueue.scala 131:10:@10597.4]
  wire  _T_10310; // @[LoadQueue.scala 131:81:@10600.4]
  wire  storesToCheck_10_15; // @[LoadQueue.scala 131:10:@10606.4]
  wire  storesToCheck_11_0; // @[LoadQueue.scala 131:10:@10648.4]
  wire  _T_10360; // @[LoadQueue.scala 131:81:@10651.4]
  wire  _T_10361; // @[LoadQueue.scala 131:72:@10652.4]
  wire  _T_10363; // @[LoadQueue.scala 132:33:@10653.4]
  wire  _T_10366; // @[LoadQueue.scala 132:41:@10655.4]
  wire  _T_10368; // @[LoadQueue.scala 132:9:@10656.4]
  wire  storesToCheck_11_1; // @[LoadQueue.scala 131:10:@10657.4]
  wire  _T_10374; // @[LoadQueue.scala 131:81:@10660.4]
  wire  _T_10375; // @[LoadQueue.scala 131:72:@10661.4]
  wire  _T_10377; // @[LoadQueue.scala 132:33:@10662.4]
  wire  _T_10380; // @[LoadQueue.scala 132:41:@10664.4]
  wire  _T_10382; // @[LoadQueue.scala 132:9:@10665.4]
  wire  storesToCheck_11_2; // @[LoadQueue.scala 131:10:@10666.4]
  wire  _T_10388; // @[LoadQueue.scala 131:81:@10669.4]
  wire  _T_10389; // @[LoadQueue.scala 131:72:@10670.4]
  wire  _T_10391; // @[LoadQueue.scala 132:33:@10671.4]
  wire  _T_10394; // @[LoadQueue.scala 132:41:@10673.4]
  wire  _T_10396; // @[LoadQueue.scala 132:9:@10674.4]
  wire  storesToCheck_11_3; // @[LoadQueue.scala 131:10:@10675.4]
  wire  _T_10402; // @[LoadQueue.scala 131:81:@10678.4]
  wire  _T_10403; // @[LoadQueue.scala 131:72:@10679.4]
  wire  _T_10405; // @[LoadQueue.scala 132:33:@10680.4]
  wire  _T_10408; // @[LoadQueue.scala 132:41:@10682.4]
  wire  _T_10410; // @[LoadQueue.scala 132:9:@10683.4]
  wire  storesToCheck_11_4; // @[LoadQueue.scala 131:10:@10684.4]
  wire  _T_10416; // @[LoadQueue.scala 131:81:@10687.4]
  wire  _T_10417; // @[LoadQueue.scala 131:72:@10688.4]
  wire  _T_10419; // @[LoadQueue.scala 132:33:@10689.4]
  wire  _T_10422; // @[LoadQueue.scala 132:41:@10691.4]
  wire  _T_10424; // @[LoadQueue.scala 132:9:@10692.4]
  wire  storesToCheck_11_5; // @[LoadQueue.scala 131:10:@10693.4]
  wire  _T_10430; // @[LoadQueue.scala 131:81:@10696.4]
  wire  _T_10431; // @[LoadQueue.scala 131:72:@10697.4]
  wire  _T_10433; // @[LoadQueue.scala 132:33:@10698.4]
  wire  _T_10436; // @[LoadQueue.scala 132:41:@10700.4]
  wire  _T_10438; // @[LoadQueue.scala 132:9:@10701.4]
  wire  storesToCheck_11_6; // @[LoadQueue.scala 131:10:@10702.4]
  wire  _T_10444; // @[LoadQueue.scala 131:81:@10705.4]
  wire  _T_10445; // @[LoadQueue.scala 131:72:@10706.4]
  wire  _T_10447; // @[LoadQueue.scala 132:33:@10707.4]
  wire  _T_10450; // @[LoadQueue.scala 132:41:@10709.4]
  wire  _T_10452; // @[LoadQueue.scala 132:9:@10710.4]
  wire  storesToCheck_11_7; // @[LoadQueue.scala 131:10:@10711.4]
  wire  _T_10458; // @[LoadQueue.scala 131:81:@10714.4]
  wire  _T_10459; // @[LoadQueue.scala 131:72:@10715.4]
  wire  _T_10461; // @[LoadQueue.scala 132:33:@10716.4]
  wire  _T_10464; // @[LoadQueue.scala 132:41:@10718.4]
  wire  _T_10466; // @[LoadQueue.scala 132:9:@10719.4]
  wire  storesToCheck_11_8; // @[LoadQueue.scala 131:10:@10720.4]
  wire  _T_10472; // @[LoadQueue.scala 131:81:@10723.4]
  wire  _T_10473; // @[LoadQueue.scala 131:72:@10724.4]
  wire  _T_10475; // @[LoadQueue.scala 132:33:@10725.4]
  wire  _T_10478; // @[LoadQueue.scala 132:41:@10727.4]
  wire  _T_10480; // @[LoadQueue.scala 132:9:@10728.4]
  wire  storesToCheck_11_9; // @[LoadQueue.scala 131:10:@10729.4]
  wire  _T_10486; // @[LoadQueue.scala 131:81:@10732.4]
  wire  _T_10487; // @[LoadQueue.scala 131:72:@10733.4]
  wire  _T_10489; // @[LoadQueue.scala 132:33:@10734.4]
  wire  _T_10492; // @[LoadQueue.scala 132:41:@10736.4]
  wire  _T_10494; // @[LoadQueue.scala 132:9:@10737.4]
  wire  storesToCheck_11_10; // @[LoadQueue.scala 131:10:@10738.4]
  wire  _T_10500; // @[LoadQueue.scala 131:81:@10741.4]
  wire  _T_10501; // @[LoadQueue.scala 131:72:@10742.4]
  wire  _T_10503; // @[LoadQueue.scala 132:33:@10743.4]
  wire  _T_10506; // @[LoadQueue.scala 132:41:@10745.4]
  wire  _T_10508; // @[LoadQueue.scala 132:9:@10746.4]
  wire  storesToCheck_11_11; // @[LoadQueue.scala 131:10:@10747.4]
  wire  _T_10514; // @[LoadQueue.scala 131:81:@10750.4]
  wire  _T_10515; // @[LoadQueue.scala 131:72:@10751.4]
  wire  _T_10517; // @[LoadQueue.scala 132:33:@10752.4]
  wire  _T_10520; // @[LoadQueue.scala 132:41:@10754.4]
  wire  _T_10522; // @[LoadQueue.scala 132:9:@10755.4]
  wire  storesToCheck_11_12; // @[LoadQueue.scala 131:10:@10756.4]
  wire  _T_10528; // @[LoadQueue.scala 131:81:@10759.4]
  wire  _T_10529; // @[LoadQueue.scala 131:72:@10760.4]
  wire  _T_10531; // @[LoadQueue.scala 132:33:@10761.4]
  wire  _T_10534; // @[LoadQueue.scala 132:41:@10763.4]
  wire  _T_10536; // @[LoadQueue.scala 132:9:@10764.4]
  wire  storesToCheck_11_13; // @[LoadQueue.scala 131:10:@10765.4]
  wire  _T_10542; // @[LoadQueue.scala 131:81:@10768.4]
  wire  _T_10543; // @[LoadQueue.scala 131:72:@10769.4]
  wire  _T_10545; // @[LoadQueue.scala 132:33:@10770.4]
  wire  _T_10548; // @[LoadQueue.scala 132:41:@10772.4]
  wire  _T_10550; // @[LoadQueue.scala 132:9:@10773.4]
  wire  storesToCheck_11_14; // @[LoadQueue.scala 131:10:@10774.4]
  wire  _T_10556; // @[LoadQueue.scala 131:81:@10777.4]
  wire  storesToCheck_11_15; // @[LoadQueue.scala 131:10:@10783.4]
  wire  storesToCheck_12_0; // @[LoadQueue.scala 131:10:@10825.4]
  wire  _T_10606; // @[LoadQueue.scala 131:81:@10828.4]
  wire  _T_10607; // @[LoadQueue.scala 131:72:@10829.4]
  wire  _T_10609; // @[LoadQueue.scala 132:33:@10830.4]
  wire  _T_10612; // @[LoadQueue.scala 132:41:@10832.4]
  wire  _T_10614; // @[LoadQueue.scala 132:9:@10833.4]
  wire  storesToCheck_12_1; // @[LoadQueue.scala 131:10:@10834.4]
  wire  _T_10620; // @[LoadQueue.scala 131:81:@10837.4]
  wire  _T_10621; // @[LoadQueue.scala 131:72:@10838.4]
  wire  _T_10623; // @[LoadQueue.scala 132:33:@10839.4]
  wire  _T_10626; // @[LoadQueue.scala 132:41:@10841.4]
  wire  _T_10628; // @[LoadQueue.scala 132:9:@10842.4]
  wire  storesToCheck_12_2; // @[LoadQueue.scala 131:10:@10843.4]
  wire  _T_10634; // @[LoadQueue.scala 131:81:@10846.4]
  wire  _T_10635; // @[LoadQueue.scala 131:72:@10847.4]
  wire  _T_10637; // @[LoadQueue.scala 132:33:@10848.4]
  wire  _T_10640; // @[LoadQueue.scala 132:41:@10850.4]
  wire  _T_10642; // @[LoadQueue.scala 132:9:@10851.4]
  wire  storesToCheck_12_3; // @[LoadQueue.scala 131:10:@10852.4]
  wire  _T_10648; // @[LoadQueue.scala 131:81:@10855.4]
  wire  _T_10649; // @[LoadQueue.scala 131:72:@10856.4]
  wire  _T_10651; // @[LoadQueue.scala 132:33:@10857.4]
  wire  _T_10654; // @[LoadQueue.scala 132:41:@10859.4]
  wire  _T_10656; // @[LoadQueue.scala 132:9:@10860.4]
  wire  storesToCheck_12_4; // @[LoadQueue.scala 131:10:@10861.4]
  wire  _T_10662; // @[LoadQueue.scala 131:81:@10864.4]
  wire  _T_10663; // @[LoadQueue.scala 131:72:@10865.4]
  wire  _T_10665; // @[LoadQueue.scala 132:33:@10866.4]
  wire  _T_10668; // @[LoadQueue.scala 132:41:@10868.4]
  wire  _T_10670; // @[LoadQueue.scala 132:9:@10869.4]
  wire  storesToCheck_12_5; // @[LoadQueue.scala 131:10:@10870.4]
  wire  _T_10676; // @[LoadQueue.scala 131:81:@10873.4]
  wire  _T_10677; // @[LoadQueue.scala 131:72:@10874.4]
  wire  _T_10679; // @[LoadQueue.scala 132:33:@10875.4]
  wire  _T_10682; // @[LoadQueue.scala 132:41:@10877.4]
  wire  _T_10684; // @[LoadQueue.scala 132:9:@10878.4]
  wire  storesToCheck_12_6; // @[LoadQueue.scala 131:10:@10879.4]
  wire  _T_10690; // @[LoadQueue.scala 131:81:@10882.4]
  wire  _T_10691; // @[LoadQueue.scala 131:72:@10883.4]
  wire  _T_10693; // @[LoadQueue.scala 132:33:@10884.4]
  wire  _T_10696; // @[LoadQueue.scala 132:41:@10886.4]
  wire  _T_10698; // @[LoadQueue.scala 132:9:@10887.4]
  wire  storesToCheck_12_7; // @[LoadQueue.scala 131:10:@10888.4]
  wire  _T_10704; // @[LoadQueue.scala 131:81:@10891.4]
  wire  _T_10705; // @[LoadQueue.scala 131:72:@10892.4]
  wire  _T_10707; // @[LoadQueue.scala 132:33:@10893.4]
  wire  _T_10710; // @[LoadQueue.scala 132:41:@10895.4]
  wire  _T_10712; // @[LoadQueue.scala 132:9:@10896.4]
  wire  storesToCheck_12_8; // @[LoadQueue.scala 131:10:@10897.4]
  wire  _T_10718; // @[LoadQueue.scala 131:81:@10900.4]
  wire  _T_10719; // @[LoadQueue.scala 131:72:@10901.4]
  wire  _T_10721; // @[LoadQueue.scala 132:33:@10902.4]
  wire  _T_10724; // @[LoadQueue.scala 132:41:@10904.4]
  wire  _T_10726; // @[LoadQueue.scala 132:9:@10905.4]
  wire  storesToCheck_12_9; // @[LoadQueue.scala 131:10:@10906.4]
  wire  _T_10732; // @[LoadQueue.scala 131:81:@10909.4]
  wire  _T_10733; // @[LoadQueue.scala 131:72:@10910.4]
  wire  _T_10735; // @[LoadQueue.scala 132:33:@10911.4]
  wire  _T_10738; // @[LoadQueue.scala 132:41:@10913.4]
  wire  _T_10740; // @[LoadQueue.scala 132:9:@10914.4]
  wire  storesToCheck_12_10; // @[LoadQueue.scala 131:10:@10915.4]
  wire  _T_10746; // @[LoadQueue.scala 131:81:@10918.4]
  wire  _T_10747; // @[LoadQueue.scala 131:72:@10919.4]
  wire  _T_10749; // @[LoadQueue.scala 132:33:@10920.4]
  wire  _T_10752; // @[LoadQueue.scala 132:41:@10922.4]
  wire  _T_10754; // @[LoadQueue.scala 132:9:@10923.4]
  wire  storesToCheck_12_11; // @[LoadQueue.scala 131:10:@10924.4]
  wire  _T_10760; // @[LoadQueue.scala 131:81:@10927.4]
  wire  _T_10761; // @[LoadQueue.scala 131:72:@10928.4]
  wire  _T_10763; // @[LoadQueue.scala 132:33:@10929.4]
  wire  _T_10766; // @[LoadQueue.scala 132:41:@10931.4]
  wire  _T_10768; // @[LoadQueue.scala 132:9:@10932.4]
  wire  storesToCheck_12_12; // @[LoadQueue.scala 131:10:@10933.4]
  wire  _T_10774; // @[LoadQueue.scala 131:81:@10936.4]
  wire  _T_10775; // @[LoadQueue.scala 131:72:@10937.4]
  wire  _T_10777; // @[LoadQueue.scala 132:33:@10938.4]
  wire  _T_10780; // @[LoadQueue.scala 132:41:@10940.4]
  wire  _T_10782; // @[LoadQueue.scala 132:9:@10941.4]
  wire  storesToCheck_12_13; // @[LoadQueue.scala 131:10:@10942.4]
  wire  _T_10788; // @[LoadQueue.scala 131:81:@10945.4]
  wire  _T_10789; // @[LoadQueue.scala 131:72:@10946.4]
  wire  _T_10791; // @[LoadQueue.scala 132:33:@10947.4]
  wire  _T_10794; // @[LoadQueue.scala 132:41:@10949.4]
  wire  _T_10796; // @[LoadQueue.scala 132:9:@10950.4]
  wire  storesToCheck_12_14; // @[LoadQueue.scala 131:10:@10951.4]
  wire  _T_10802; // @[LoadQueue.scala 131:81:@10954.4]
  wire  storesToCheck_12_15; // @[LoadQueue.scala 131:10:@10960.4]
  wire  storesToCheck_13_0; // @[LoadQueue.scala 131:10:@11002.4]
  wire  _T_10852; // @[LoadQueue.scala 131:81:@11005.4]
  wire  _T_10853; // @[LoadQueue.scala 131:72:@11006.4]
  wire  _T_10855; // @[LoadQueue.scala 132:33:@11007.4]
  wire  _T_10858; // @[LoadQueue.scala 132:41:@11009.4]
  wire  _T_10860; // @[LoadQueue.scala 132:9:@11010.4]
  wire  storesToCheck_13_1; // @[LoadQueue.scala 131:10:@11011.4]
  wire  _T_10866; // @[LoadQueue.scala 131:81:@11014.4]
  wire  _T_10867; // @[LoadQueue.scala 131:72:@11015.4]
  wire  _T_10869; // @[LoadQueue.scala 132:33:@11016.4]
  wire  _T_10872; // @[LoadQueue.scala 132:41:@11018.4]
  wire  _T_10874; // @[LoadQueue.scala 132:9:@11019.4]
  wire  storesToCheck_13_2; // @[LoadQueue.scala 131:10:@11020.4]
  wire  _T_10880; // @[LoadQueue.scala 131:81:@11023.4]
  wire  _T_10881; // @[LoadQueue.scala 131:72:@11024.4]
  wire  _T_10883; // @[LoadQueue.scala 132:33:@11025.4]
  wire  _T_10886; // @[LoadQueue.scala 132:41:@11027.4]
  wire  _T_10888; // @[LoadQueue.scala 132:9:@11028.4]
  wire  storesToCheck_13_3; // @[LoadQueue.scala 131:10:@11029.4]
  wire  _T_10894; // @[LoadQueue.scala 131:81:@11032.4]
  wire  _T_10895; // @[LoadQueue.scala 131:72:@11033.4]
  wire  _T_10897; // @[LoadQueue.scala 132:33:@11034.4]
  wire  _T_10900; // @[LoadQueue.scala 132:41:@11036.4]
  wire  _T_10902; // @[LoadQueue.scala 132:9:@11037.4]
  wire  storesToCheck_13_4; // @[LoadQueue.scala 131:10:@11038.4]
  wire  _T_10908; // @[LoadQueue.scala 131:81:@11041.4]
  wire  _T_10909; // @[LoadQueue.scala 131:72:@11042.4]
  wire  _T_10911; // @[LoadQueue.scala 132:33:@11043.4]
  wire  _T_10914; // @[LoadQueue.scala 132:41:@11045.4]
  wire  _T_10916; // @[LoadQueue.scala 132:9:@11046.4]
  wire  storesToCheck_13_5; // @[LoadQueue.scala 131:10:@11047.4]
  wire  _T_10922; // @[LoadQueue.scala 131:81:@11050.4]
  wire  _T_10923; // @[LoadQueue.scala 131:72:@11051.4]
  wire  _T_10925; // @[LoadQueue.scala 132:33:@11052.4]
  wire  _T_10928; // @[LoadQueue.scala 132:41:@11054.4]
  wire  _T_10930; // @[LoadQueue.scala 132:9:@11055.4]
  wire  storesToCheck_13_6; // @[LoadQueue.scala 131:10:@11056.4]
  wire  _T_10936; // @[LoadQueue.scala 131:81:@11059.4]
  wire  _T_10937; // @[LoadQueue.scala 131:72:@11060.4]
  wire  _T_10939; // @[LoadQueue.scala 132:33:@11061.4]
  wire  _T_10942; // @[LoadQueue.scala 132:41:@11063.4]
  wire  _T_10944; // @[LoadQueue.scala 132:9:@11064.4]
  wire  storesToCheck_13_7; // @[LoadQueue.scala 131:10:@11065.4]
  wire  _T_10950; // @[LoadQueue.scala 131:81:@11068.4]
  wire  _T_10951; // @[LoadQueue.scala 131:72:@11069.4]
  wire  _T_10953; // @[LoadQueue.scala 132:33:@11070.4]
  wire  _T_10956; // @[LoadQueue.scala 132:41:@11072.4]
  wire  _T_10958; // @[LoadQueue.scala 132:9:@11073.4]
  wire  storesToCheck_13_8; // @[LoadQueue.scala 131:10:@11074.4]
  wire  _T_10964; // @[LoadQueue.scala 131:81:@11077.4]
  wire  _T_10965; // @[LoadQueue.scala 131:72:@11078.4]
  wire  _T_10967; // @[LoadQueue.scala 132:33:@11079.4]
  wire  _T_10970; // @[LoadQueue.scala 132:41:@11081.4]
  wire  _T_10972; // @[LoadQueue.scala 132:9:@11082.4]
  wire  storesToCheck_13_9; // @[LoadQueue.scala 131:10:@11083.4]
  wire  _T_10978; // @[LoadQueue.scala 131:81:@11086.4]
  wire  _T_10979; // @[LoadQueue.scala 131:72:@11087.4]
  wire  _T_10981; // @[LoadQueue.scala 132:33:@11088.4]
  wire  _T_10984; // @[LoadQueue.scala 132:41:@11090.4]
  wire  _T_10986; // @[LoadQueue.scala 132:9:@11091.4]
  wire  storesToCheck_13_10; // @[LoadQueue.scala 131:10:@11092.4]
  wire  _T_10992; // @[LoadQueue.scala 131:81:@11095.4]
  wire  _T_10993; // @[LoadQueue.scala 131:72:@11096.4]
  wire  _T_10995; // @[LoadQueue.scala 132:33:@11097.4]
  wire  _T_10998; // @[LoadQueue.scala 132:41:@11099.4]
  wire  _T_11000; // @[LoadQueue.scala 132:9:@11100.4]
  wire  storesToCheck_13_11; // @[LoadQueue.scala 131:10:@11101.4]
  wire  _T_11006; // @[LoadQueue.scala 131:81:@11104.4]
  wire  _T_11007; // @[LoadQueue.scala 131:72:@11105.4]
  wire  _T_11009; // @[LoadQueue.scala 132:33:@11106.4]
  wire  _T_11012; // @[LoadQueue.scala 132:41:@11108.4]
  wire  _T_11014; // @[LoadQueue.scala 132:9:@11109.4]
  wire  storesToCheck_13_12; // @[LoadQueue.scala 131:10:@11110.4]
  wire  _T_11020; // @[LoadQueue.scala 131:81:@11113.4]
  wire  _T_11021; // @[LoadQueue.scala 131:72:@11114.4]
  wire  _T_11023; // @[LoadQueue.scala 132:33:@11115.4]
  wire  _T_11026; // @[LoadQueue.scala 132:41:@11117.4]
  wire  _T_11028; // @[LoadQueue.scala 132:9:@11118.4]
  wire  storesToCheck_13_13; // @[LoadQueue.scala 131:10:@11119.4]
  wire  _T_11034; // @[LoadQueue.scala 131:81:@11122.4]
  wire  _T_11035; // @[LoadQueue.scala 131:72:@11123.4]
  wire  _T_11037; // @[LoadQueue.scala 132:33:@11124.4]
  wire  _T_11040; // @[LoadQueue.scala 132:41:@11126.4]
  wire  _T_11042; // @[LoadQueue.scala 132:9:@11127.4]
  wire  storesToCheck_13_14; // @[LoadQueue.scala 131:10:@11128.4]
  wire  _T_11048; // @[LoadQueue.scala 131:81:@11131.4]
  wire  storesToCheck_13_15; // @[LoadQueue.scala 131:10:@11137.4]
  wire  storesToCheck_14_0; // @[LoadQueue.scala 131:10:@11179.4]
  wire  _T_11098; // @[LoadQueue.scala 131:81:@11182.4]
  wire  _T_11099; // @[LoadQueue.scala 131:72:@11183.4]
  wire  _T_11101; // @[LoadQueue.scala 132:33:@11184.4]
  wire  _T_11104; // @[LoadQueue.scala 132:41:@11186.4]
  wire  _T_11106; // @[LoadQueue.scala 132:9:@11187.4]
  wire  storesToCheck_14_1; // @[LoadQueue.scala 131:10:@11188.4]
  wire  _T_11112; // @[LoadQueue.scala 131:81:@11191.4]
  wire  _T_11113; // @[LoadQueue.scala 131:72:@11192.4]
  wire  _T_11115; // @[LoadQueue.scala 132:33:@11193.4]
  wire  _T_11118; // @[LoadQueue.scala 132:41:@11195.4]
  wire  _T_11120; // @[LoadQueue.scala 132:9:@11196.4]
  wire  storesToCheck_14_2; // @[LoadQueue.scala 131:10:@11197.4]
  wire  _T_11126; // @[LoadQueue.scala 131:81:@11200.4]
  wire  _T_11127; // @[LoadQueue.scala 131:72:@11201.4]
  wire  _T_11129; // @[LoadQueue.scala 132:33:@11202.4]
  wire  _T_11132; // @[LoadQueue.scala 132:41:@11204.4]
  wire  _T_11134; // @[LoadQueue.scala 132:9:@11205.4]
  wire  storesToCheck_14_3; // @[LoadQueue.scala 131:10:@11206.4]
  wire  _T_11140; // @[LoadQueue.scala 131:81:@11209.4]
  wire  _T_11141; // @[LoadQueue.scala 131:72:@11210.4]
  wire  _T_11143; // @[LoadQueue.scala 132:33:@11211.4]
  wire  _T_11146; // @[LoadQueue.scala 132:41:@11213.4]
  wire  _T_11148; // @[LoadQueue.scala 132:9:@11214.4]
  wire  storesToCheck_14_4; // @[LoadQueue.scala 131:10:@11215.4]
  wire  _T_11154; // @[LoadQueue.scala 131:81:@11218.4]
  wire  _T_11155; // @[LoadQueue.scala 131:72:@11219.4]
  wire  _T_11157; // @[LoadQueue.scala 132:33:@11220.4]
  wire  _T_11160; // @[LoadQueue.scala 132:41:@11222.4]
  wire  _T_11162; // @[LoadQueue.scala 132:9:@11223.4]
  wire  storesToCheck_14_5; // @[LoadQueue.scala 131:10:@11224.4]
  wire  _T_11168; // @[LoadQueue.scala 131:81:@11227.4]
  wire  _T_11169; // @[LoadQueue.scala 131:72:@11228.4]
  wire  _T_11171; // @[LoadQueue.scala 132:33:@11229.4]
  wire  _T_11174; // @[LoadQueue.scala 132:41:@11231.4]
  wire  _T_11176; // @[LoadQueue.scala 132:9:@11232.4]
  wire  storesToCheck_14_6; // @[LoadQueue.scala 131:10:@11233.4]
  wire  _T_11182; // @[LoadQueue.scala 131:81:@11236.4]
  wire  _T_11183; // @[LoadQueue.scala 131:72:@11237.4]
  wire  _T_11185; // @[LoadQueue.scala 132:33:@11238.4]
  wire  _T_11188; // @[LoadQueue.scala 132:41:@11240.4]
  wire  _T_11190; // @[LoadQueue.scala 132:9:@11241.4]
  wire  storesToCheck_14_7; // @[LoadQueue.scala 131:10:@11242.4]
  wire  _T_11196; // @[LoadQueue.scala 131:81:@11245.4]
  wire  _T_11197; // @[LoadQueue.scala 131:72:@11246.4]
  wire  _T_11199; // @[LoadQueue.scala 132:33:@11247.4]
  wire  _T_11202; // @[LoadQueue.scala 132:41:@11249.4]
  wire  _T_11204; // @[LoadQueue.scala 132:9:@11250.4]
  wire  storesToCheck_14_8; // @[LoadQueue.scala 131:10:@11251.4]
  wire  _T_11210; // @[LoadQueue.scala 131:81:@11254.4]
  wire  _T_11211; // @[LoadQueue.scala 131:72:@11255.4]
  wire  _T_11213; // @[LoadQueue.scala 132:33:@11256.4]
  wire  _T_11216; // @[LoadQueue.scala 132:41:@11258.4]
  wire  _T_11218; // @[LoadQueue.scala 132:9:@11259.4]
  wire  storesToCheck_14_9; // @[LoadQueue.scala 131:10:@11260.4]
  wire  _T_11224; // @[LoadQueue.scala 131:81:@11263.4]
  wire  _T_11225; // @[LoadQueue.scala 131:72:@11264.4]
  wire  _T_11227; // @[LoadQueue.scala 132:33:@11265.4]
  wire  _T_11230; // @[LoadQueue.scala 132:41:@11267.4]
  wire  _T_11232; // @[LoadQueue.scala 132:9:@11268.4]
  wire  storesToCheck_14_10; // @[LoadQueue.scala 131:10:@11269.4]
  wire  _T_11238; // @[LoadQueue.scala 131:81:@11272.4]
  wire  _T_11239; // @[LoadQueue.scala 131:72:@11273.4]
  wire  _T_11241; // @[LoadQueue.scala 132:33:@11274.4]
  wire  _T_11244; // @[LoadQueue.scala 132:41:@11276.4]
  wire  _T_11246; // @[LoadQueue.scala 132:9:@11277.4]
  wire  storesToCheck_14_11; // @[LoadQueue.scala 131:10:@11278.4]
  wire  _T_11252; // @[LoadQueue.scala 131:81:@11281.4]
  wire  _T_11253; // @[LoadQueue.scala 131:72:@11282.4]
  wire  _T_11255; // @[LoadQueue.scala 132:33:@11283.4]
  wire  _T_11258; // @[LoadQueue.scala 132:41:@11285.4]
  wire  _T_11260; // @[LoadQueue.scala 132:9:@11286.4]
  wire  storesToCheck_14_12; // @[LoadQueue.scala 131:10:@11287.4]
  wire  _T_11266; // @[LoadQueue.scala 131:81:@11290.4]
  wire  _T_11267; // @[LoadQueue.scala 131:72:@11291.4]
  wire  _T_11269; // @[LoadQueue.scala 132:33:@11292.4]
  wire  _T_11272; // @[LoadQueue.scala 132:41:@11294.4]
  wire  _T_11274; // @[LoadQueue.scala 132:9:@11295.4]
  wire  storesToCheck_14_13; // @[LoadQueue.scala 131:10:@11296.4]
  wire  _T_11280; // @[LoadQueue.scala 131:81:@11299.4]
  wire  _T_11281; // @[LoadQueue.scala 131:72:@11300.4]
  wire  _T_11283; // @[LoadQueue.scala 132:33:@11301.4]
  wire  _T_11286; // @[LoadQueue.scala 132:41:@11303.4]
  wire  _T_11288; // @[LoadQueue.scala 132:9:@11304.4]
  wire  storesToCheck_14_14; // @[LoadQueue.scala 131:10:@11305.4]
  wire  _T_11294; // @[LoadQueue.scala 131:81:@11308.4]
  wire  storesToCheck_14_15; // @[LoadQueue.scala 131:10:@11314.4]
  wire  storesToCheck_15_0; // @[LoadQueue.scala 131:10:@11356.4]
  wire  _T_11344; // @[LoadQueue.scala 131:81:@11359.4]
  wire  _T_11345; // @[LoadQueue.scala 131:72:@11360.4]
  wire  _T_11347; // @[LoadQueue.scala 132:33:@11361.4]
  wire  _T_11350; // @[LoadQueue.scala 132:41:@11363.4]
  wire  _T_11352; // @[LoadQueue.scala 132:9:@11364.4]
  wire  storesToCheck_15_1; // @[LoadQueue.scala 131:10:@11365.4]
  wire  _T_11358; // @[LoadQueue.scala 131:81:@11368.4]
  wire  _T_11359; // @[LoadQueue.scala 131:72:@11369.4]
  wire  _T_11361; // @[LoadQueue.scala 132:33:@11370.4]
  wire  _T_11364; // @[LoadQueue.scala 132:41:@11372.4]
  wire  _T_11366; // @[LoadQueue.scala 132:9:@11373.4]
  wire  storesToCheck_15_2; // @[LoadQueue.scala 131:10:@11374.4]
  wire  _T_11372; // @[LoadQueue.scala 131:81:@11377.4]
  wire  _T_11373; // @[LoadQueue.scala 131:72:@11378.4]
  wire  _T_11375; // @[LoadQueue.scala 132:33:@11379.4]
  wire  _T_11378; // @[LoadQueue.scala 132:41:@11381.4]
  wire  _T_11380; // @[LoadQueue.scala 132:9:@11382.4]
  wire  storesToCheck_15_3; // @[LoadQueue.scala 131:10:@11383.4]
  wire  _T_11386; // @[LoadQueue.scala 131:81:@11386.4]
  wire  _T_11387; // @[LoadQueue.scala 131:72:@11387.4]
  wire  _T_11389; // @[LoadQueue.scala 132:33:@11388.4]
  wire  _T_11392; // @[LoadQueue.scala 132:41:@11390.4]
  wire  _T_11394; // @[LoadQueue.scala 132:9:@11391.4]
  wire  storesToCheck_15_4; // @[LoadQueue.scala 131:10:@11392.4]
  wire  _T_11400; // @[LoadQueue.scala 131:81:@11395.4]
  wire  _T_11401; // @[LoadQueue.scala 131:72:@11396.4]
  wire  _T_11403; // @[LoadQueue.scala 132:33:@11397.4]
  wire  _T_11406; // @[LoadQueue.scala 132:41:@11399.4]
  wire  _T_11408; // @[LoadQueue.scala 132:9:@11400.4]
  wire  storesToCheck_15_5; // @[LoadQueue.scala 131:10:@11401.4]
  wire  _T_11414; // @[LoadQueue.scala 131:81:@11404.4]
  wire  _T_11415; // @[LoadQueue.scala 131:72:@11405.4]
  wire  _T_11417; // @[LoadQueue.scala 132:33:@11406.4]
  wire  _T_11420; // @[LoadQueue.scala 132:41:@11408.4]
  wire  _T_11422; // @[LoadQueue.scala 132:9:@11409.4]
  wire  storesToCheck_15_6; // @[LoadQueue.scala 131:10:@11410.4]
  wire  _T_11428; // @[LoadQueue.scala 131:81:@11413.4]
  wire  _T_11429; // @[LoadQueue.scala 131:72:@11414.4]
  wire  _T_11431; // @[LoadQueue.scala 132:33:@11415.4]
  wire  _T_11434; // @[LoadQueue.scala 132:41:@11417.4]
  wire  _T_11436; // @[LoadQueue.scala 132:9:@11418.4]
  wire  storesToCheck_15_7; // @[LoadQueue.scala 131:10:@11419.4]
  wire  _T_11442; // @[LoadQueue.scala 131:81:@11422.4]
  wire  _T_11443; // @[LoadQueue.scala 131:72:@11423.4]
  wire  _T_11445; // @[LoadQueue.scala 132:33:@11424.4]
  wire  _T_11448; // @[LoadQueue.scala 132:41:@11426.4]
  wire  _T_11450; // @[LoadQueue.scala 132:9:@11427.4]
  wire  storesToCheck_15_8; // @[LoadQueue.scala 131:10:@11428.4]
  wire  _T_11456; // @[LoadQueue.scala 131:81:@11431.4]
  wire  _T_11457; // @[LoadQueue.scala 131:72:@11432.4]
  wire  _T_11459; // @[LoadQueue.scala 132:33:@11433.4]
  wire  _T_11462; // @[LoadQueue.scala 132:41:@11435.4]
  wire  _T_11464; // @[LoadQueue.scala 132:9:@11436.4]
  wire  storesToCheck_15_9; // @[LoadQueue.scala 131:10:@11437.4]
  wire  _T_11470; // @[LoadQueue.scala 131:81:@11440.4]
  wire  _T_11471; // @[LoadQueue.scala 131:72:@11441.4]
  wire  _T_11473; // @[LoadQueue.scala 132:33:@11442.4]
  wire  _T_11476; // @[LoadQueue.scala 132:41:@11444.4]
  wire  _T_11478; // @[LoadQueue.scala 132:9:@11445.4]
  wire  storesToCheck_15_10; // @[LoadQueue.scala 131:10:@11446.4]
  wire  _T_11484; // @[LoadQueue.scala 131:81:@11449.4]
  wire  _T_11485; // @[LoadQueue.scala 131:72:@11450.4]
  wire  _T_11487; // @[LoadQueue.scala 132:33:@11451.4]
  wire  _T_11490; // @[LoadQueue.scala 132:41:@11453.4]
  wire  _T_11492; // @[LoadQueue.scala 132:9:@11454.4]
  wire  storesToCheck_15_11; // @[LoadQueue.scala 131:10:@11455.4]
  wire  _T_11498; // @[LoadQueue.scala 131:81:@11458.4]
  wire  _T_11499; // @[LoadQueue.scala 131:72:@11459.4]
  wire  _T_11501; // @[LoadQueue.scala 132:33:@11460.4]
  wire  _T_11504; // @[LoadQueue.scala 132:41:@11462.4]
  wire  _T_11506; // @[LoadQueue.scala 132:9:@11463.4]
  wire  storesToCheck_15_12; // @[LoadQueue.scala 131:10:@11464.4]
  wire  _T_11512; // @[LoadQueue.scala 131:81:@11467.4]
  wire  _T_11513; // @[LoadQueue.scala 131:72:@11468.4]
  wire  _T_11515; // @[LoadQueue.scala 132:33:@11469.4]
  wire  _T_11518; // @[LoadQueue.scala 132:41:@11471.4]
  wire  _T_11520; // @[LoadQueue.scala 132:9:@11472.4]
  wire  storesToCheck_15_13; // @[LoadQueue.scala 131:10:@11473.4]
  wire  _T_11526; // @[LoadQueue.scala 131:81:@11476.4]
  wire  _T_11527; // @[LoadQueue.scala 131:72:@11477.4]
  wire  _T_11529; // @[LoadQueue.scala 132:33:@11478.4]
  wire  _T_11532; // @[LoadQueue.scala 132:41:@11480.4]
  wire  _T_11534; // @[LoadQueue.scala 132:9:@11481.4]
  wire  storesToCheck_15_14; // @[LoadQueue.scala 131:10:@11482.4]
  wire  _T_11540; // @[LoadQueue.scala 131:81:@11485.4]
  wire  storesToCheck_15_15; // @[LoadQueue.scala 131:10:@11491.4]
  wire  _T_12802; // @[LoadQueue.scala 141:18:@11526.4]
  wire  entriesToCheck_0_0; // @[LoadQueue.scala 141:26:@11527.4]
  wire  _T_12804; // @[LoadQueue.scala 141:18:@11528.4]
  wire  entriesToCheck_0_1; // @[LoadQueue.scala 141:26:@11529.4]
  wire  _T_12806; // @[LoadQueue.scala 141:18:@11530.4]
  wire  entriesToCheck_0_2; // @[LoadQueue.scala 141:26:@11531.4]
  wire  _T_12808; // @[LoadQueue.scala 141:18:@11532.4]
  wire  entriesToCheck_0_3; // @[LoadQueue.scala 141:26:@11533.4]
  wire  _T_12810; // @[LoadQueue.scala 141:18:@11534.4]
  wire  entriesToCheck_0_4; // @[LoadQueue.scala 141:26:@11535.4]
  wire  _T_12812; // @[LoadQueue.scala 141:18:@11536.4]
  wire  entriesToCheck_0_5; // @[LoadQueue.scala 141:26:@11537.4]
  wire  _T_12814; // @[LoadQueue.scala 141:18:@11538.4]
  wire  entriesToCheck_0_6; // @[LoadQueue.scala 141:26:@11539.4]
  wire  _T_12816; // @[LoadQueue.scala 141:18:@11540.4]
  wire  entriesToCheck_0_7; // @[LoadQueue.scala 141:26:@11541.4]
  wire  _T_12818; // @[LoadQueue.scala 141:18:@11542.4]
  wire  entriesToCheck_0_8; // @[LoadQueue.scala 141:26:@11543.4]
  wire  _T_12820; // @[LoadQueue.scala 141:18:@11544.4]
  wire  entriesToCheck_0_9; // @[LoadQueue.scala 141:26:@11545.4]
  wire  _T_12822; // @[LoadQueue.scala 141:18:@11546.4]
  wire  entriesToCheck_0_10; // @[LoadQueue.scala 141:26:@11547.4]
  wire  _T_12824; // @[LoadQueue.scala 141:18:@11548.4]
  wire  entriesToCheck_0_11; // @[LoadQueue.scala 141:26:@11549.4]
  wire  _T_12826; // @[LoadQueue.scala 141:18:@11550.4]
  wire  entriesToCheck_0_12; // @[LoadQueue.scala 141:26:@11551.4]
  wire  _T_12828; // @[LoadQueue.scala 141:18:@11552.4]
  wire  entriesToCheck_0_13; // @[LoadQueue.scala 141:26:@11553.4]
  wire  _T_12830; // @[LoadQueue.scala 141:18:@11554.4]
  wire  entriesToCheck_0_14; // @[LoadQueue.scala 141:26:@11555.4]
  wire  _T_12832; // @[LoadQueue.scala 141:18:@11556.4]
  wire  entriesToCheck_0_15; // @[LoadQueue.scala 141:26:@11557.4]
  wire  _T_12834; // @[LoadQueue.scala 141:18:@11574.4]
  wire  entriesToCheck_1_0; // @[LoadQueue.scala 141:26:@11575.4]
  wire  _T_12836; // @[LoadQueue.scala 141:18:@11576.4]
  wire  entriesToCheck_1_1; // @[LoadQueue.scala 141:26:@11577.4]
  wire  _T_12838; // @[LoadQueue.scala 141:18:@11578.4]
  wire  entriesToCheck_1_2; // @[LoadQueue.scala 141:26:@11579.4]
  wire  _T_12840; // @[LoadQueue.scala 141:18:@11580.4]
  wire  entriesToCheck_1_3; // @[LoadQueue.scala 141:26:@11581.4]
  wire  _T_12842; // @[LoadQueue.scala 141:18:@11582.4]
  wire  entriesToCheck_1_4; // @[LoadQueue.scala 141:26:@11583.4]
  wire  _T_12844; // @[LoadQueue.scala 141:18:@11584.4]
  wire  entriesToCheck_1_5; // @[LoadQueue.scala 141:26:@11585.4]
  wire  _T_12846; // @[LoadQueue.scala 141:18:@11586.4]
  wire  entriesToCheck_1_6; // @[LoadQueue.scala 141:26:@11587.4]
  wire  _T_12848; // @[LoadQueue.scala 141:18:@11588.4]
  wire  entriesToCheck_1_7; // @[LoadQueue.scala 141:26:@11589.4]
  wire  _T_12850; // @[LoadQueue.scala 141:18:@11590.4]
  wire  entriesToCheck_1_8; // @[LoadQueue.scala 141:26:@11591.4]
  wire  _T_12852; // @[LoadQueue.scala 141:18:@11592.4]
  wire  entriesToCheck_1_9; // @[LoadQueue.scala 141:26:@11593.4]
  wire  _T_12854; // @[LoadQueue.scala 141:18:@11594.4]
  wire  entriesToCheck_1_10; // @[LoadQueue.scala 141:26:@11595.4]
  wire  _T_12856; // @[LoadQueue.scala 141:18:@11596.4]
  wire  entriesToCheck_1_11; // @[LoadQueue.scala 141:26:@11597.4]
  wire  _T_12858; // @[LoadQueue.scala 141:18:@11598.4]
  wire  entriesToCheck_1_12; // @[LoadQueue.scala 141:26:@11599.4]
  wire  _T_12860; // @[LoadQueue.scala 141:18:@11600.4]
  wire  entriesToCheck_1_13; // @[LoadQueue.scala 141:26:@11601.4]
  wire  _T_12862; // @[LoadQueue.scala 141:18:@11602.4]
  wire  entriesToCheck_1_14; // @[LoadQueue.scala 141:26:@11603.4]
  wire  _T_12864; // @[LoadQueue.scala 141:18:@11604.4]
  wire  entriesToCheck_1_15; // @[LoadQueue.scala 141:26:@11605.4]
  wire  _T_12866; // @[LoadQueue.scala 141:18:@11622.4]
  wire  entriesToCheck_2_0; // @[LoadQueue.scala 141:26:@11623.4]
  wire  _T_12868; // @[LoadQueue.scala 141:18:@11624.4]
  wire  entriesToCheck_2_1; // @[LoadQueue.scala 141:26:@11625.4]
  wire  _T_12870; // @[LoadQueue.scala 141:18:@11626.4]
  wire  entriesToCheck_2_2; // @[LoadQueue.scala 141:26:@11627.4]
  wire  _T_12872; // @[LoadQueue.scala 141:18:@11628.4]
  wire  entriesToCheck_2_3; // @[LoadQueue.scala 141:26:@11629.4]
  wire  _T_12874; // @[LoadQueue.scala 141:18:@11630.4]
  wire  entriesToCheck_2_4; // @[LoadQueue.scala 141:26:@11631.4]
  wire  _T_12876; // @[LoadQueue.scala 141:18:@11632.4]
  wire  entriesToCheck_2_5; // @[LoadQueue.scala 141:26:@11633.4]
  wire  _T_12878; // @[LoadQueue.scala 141:18:@11634.4]
  wire  entriesToCheck_2_6; // @[LoadQueue.scala 141:26:@11635.4]
  wire  _T_12880; // @[LoadQueue.scala 141:18:@11636.4]
  wire  entriesToCheck_2_7; // @[LoadQueue.scala 141:26:@11637.4]
  wire  _T_12882; // @[LoadQueue.scala 141:18:@11638.4]
  wire  entriesToCheck_2_8; // @[LoadQueue.scala 141:26:@11639.4]
  wire  _T_12884; // @[LoadQueue.scala 141:18:@11640.4]
  wire  entriesToCheck_2_9; // @[LoadQueue.scala 141:26:@11641.4]
  wire  _T_12886; // @[LoadQueue.scala 141:18:@11642.4]
  wire  entriesToCheck_2_10; // @[LoadQueue.scala 141:26:@11643.4]
  wire  _T_12888; // @[LoadQueue.scala 141:18:@11644.4]
  wire  entriesToCheck_2_11; // @[LoadQueue.scala 141:26:@11645.4]
  wire  _T_12890; // @[LoadQueue.scala 141:18:@11646.4]
  wire  entriesToCheck_2_12; // @[LoadQueue.scala 141:26:@11647.4]
  wire  _T_12892; // @[LoadQueue.scala 141:18:@11648.4]
  wire  entriesToCheck_2_13; // @[LoadQueue.scala 141:26:@11649.4]
  wire  _T_12894; // @[LoadQueue.scala 141:18:@11650.4]
  wire  entriesToCheck_2_14; // @[LoadQueue.scala 141:26:@11651.4]
  wire  _T_12896; // @[LoadQueue.scala 141:18:@11652.4]
  wire  entriesToCheck_2_15; // @[LoadQueue.scala 141:26:@11653.4]
  wire  _T_12898; // @[LoadQueue.scala 141:18:@11670.4]
  wire  entriesToCheck_3_0; // @[LoadQueue.scala 141:26:@11671.4]
  wire  _T_12900; // @[LoadQueue.scala 141:18:@11672.4]
  wire  entriesToCheck_3_1; // @[LoadQueue.scala 141:26:@11673.4]
  wire  _T_12902; // @[LoadQueue.scala 141:18:@11674.4]
  wire  entriesToCheck_3_2; // @[LoadQueue.scala 141:26:@11675.4]
  wire  _T_12904; // @[LoadQueue.scala 141:18:@11676.4]
  wire  entriesToCheck_3_3; // @[LoadQueue.scala 141:26:@11677.4]
  wire  _T_12906; // @[LoadQueue.scala 141:18:@11678.4]
  wire  entriesToCheck_3_4; // @[LoadQueue.scala 141:26:@11679.4]
  wire  _T_12908; // @[LoadQueue.scala 141:18:@11680.4]
  wire  entriesToCheck_3_5; // @[LoadQueue.scala 141:26:@11681.4]
  wire  _T_12910; // @[LoadQueue.scala 141:18:@11682.4]
  wire  entriesToCheck_3_6; // @[LoadQueue.scala 141:26:@11683.4]
  wire  _T_12912; // @[LoadQueue.scala 141:18:@11684.4]
  wire  entriesToCheck_3_7; // @[LoadQueue.scala 141:26:@11685.4]
  wire  _T_12914; // @[LoadQueue.scala 141:18:@11686.4]
  wire  entriesToCheck_3_8; // @[LoadQueue.scala 141:26:@11687.4]
  wire  _T_12916; // @[LoadQueue.scala 141:18:@11688.4]
  wire  entriesToCheck_3_9; // @[LoadQueue.scala 141:26:@11689.4]
  wire  _T_12918; // @[LoadQueue.scala 141:18:@11690.4]
  wire  entriesToCheck_3_10; // @[LoadQueue.scala 141:26:@11691.4]
  wire  _T_12920; // @[LoadQueue.scala 141:18:@11692.4]
  wire  entriesToCheck_3_11; // @[LoadQueue.scala 141:26:@11693.4]
  wire  _T_12922; // @[LoadQueue.scala 141:18:@11694.4]
  wire  entriesToCheck_3_12; // @[LoadQueue.scala 141:26:@11695.4]
  wire  _T_12924; // @[LoadQueue.scala 141:18:@11696.4]
  wire  entriesToCheck_3_13; // @[LoadQueue.scala 141:26:@11697.4]
  wire  _T_12926; // @[LoadQueue.scala 141:18:@11698.4]
  wire  entriesToCheck_3_14; // @[LoadQueue.scala 141:26:@11699.4]
  wire  _T_12928; // @[LoadQueue.scala 141:18:@11700.4]
  wire  entriesToCheck_3_15; // @[LoadQueue.scala 141:26:@11701.4]
  wire  _T_12930; // @[LoadQueue.scala 141:18:@11718.4]
  wire  entriesToCheck_4_0; // @[LoadQueue.scala 141:26:@11719.4]
  wire  _T_12932; // @[LoadQueue.scala 141:18:@11720.4]
  wire  entriesToCheck_4_1; // @[LoadQueue.scala 141:26:@11721.4]
  wire  _T_12934; // @[LoadQueue.scala 141:18:@11722.4]
  wire  entriesToCheck_4_2; // @[LoadQueue.scala 141:26:@11723.4]
  wire  _T_12936; // @[LoadQueue.scala 141:18:@11724.4]
  wire  entriesToCheck_4_3; // @[LoadQueue.scala 141:26:@11725.4]
  wire  _T_12938; // @[LoadQueue.scala 141:18:@11726.4]
  wire  entriesToCheck_4_4; // @[LoadQueue.scala 141:26:@11727.4]
  wire  _T_12940; // @[LoadQueue.scala 141:18:@11728.4]
  wire  entriesToCheck_4_5; // @[LoadQueue.scala 141:26:@11729.4]
  wire  _T_12942; // @[LoadQueue.scala 141:18:@11730.4]
  wire  entriesToCheck_4_6; // @[LoadQueue.scala 141:26:@11731.4]
  wire  _T_12944; // @[LoadQueue.scala 141:18:@11732.4]
  wire  entriesToCheck_4_7; // @[LoadQueue.scala 141:26:@11733.4]
  wire  _T_12946; // @[LoadQueue.scala 141:18:@11734.4]
  wire  entriesToCheck_4_8; // @[LoadQueue.scala 141:26:@11735.4]
  wire  _T_12948; // @[LoadQueue.scala 141:18:@11736.4]
  wire  entriesToCheck_4_9; // @[LoadQueue.scala 141:26:@11737.4]
  wire  _T_12950; // @[LoadQueue.scala 141:18:@11738.4]
  wire  entriesToCheck_4_10; // @[LoadQueue.scala 141:26:@11739.4]
  wire  _T_12952; // @[LoadQueue.scala 141:18:@11740.4]
  wire  entriesToCheck_4_11; // @[LoadQueue.scala 141:26:@11741.4]
  wire  _T_12954; // @[LoadQueue.scala 141:18:@11742.4]
  wire  entriesToCheck_4_12; // @[LoadQueue.scala 141:26:@11743.4]
  wire  _T_12956; // @[LoadQueue.scala 141:18:@11744.4]
  wire  entriesToCheck_4_13; // @[LoadQueue.scala 141:26:@11745.4]
  wire  _T_12958; // @[LoadQueue.scala 141:18:@11746.4]
  wire  entriesToCheck_4_14; // @[LoadQueue.scala 141:26:@11747.4]
  wire  _T_12960; // @[LoadQueue.scala 141:18:@11748.4]
  wire  entriesToCheck_4_15; // @[LoadQueue.scala 141:26:@11749.4]
  wire  _T_12962; // @[LoadQueue.scala 141:18:@11766.4]
  wire  entriesToCheck_5_0; // @[LoadQueue.scala 141:26:@11767.4]
  wire  _T_12964; // @[LoadQueue.scala 141:18:@11768.4]
  wire  entriesToCheck_5_1; // @[LoadQueue.scala 141:26:@11769.4]
  wire  _T_12966; // @[LoadQueue.scala 141:18:@11770.4]
  wire  entriesToCheck_5_2; // @[LoadQueue.scala 141:26:@11771.4]
  wire  _T_12968; // @[LoadQueue.scala 141:18:@11772.4]
  wire  entriesToCheck_5_3; // @[LoadQueue.scala 141:26:@11773.4]
  wire  _T_12970; // @[LoadQueue.scala 141:18:@11774.4]
  wire  entriesToCheck_5_4; // @[LoadQueue.scala 141:26:@11775.4]
  wire  _T_12972; // @[LoadQueue.scala 141:18:@11776.4]
  wire  entriesToCheck_5_5; // @[LoadQueue.scala 141:26:@11777.4]
  wire  _T_12974; // @[LoadQueue.scala 141:18:@11778.4]
  wire  entriesToCheck_5_6; // @[LoadQueue.scala 141:26:@11779.4]
  wire  _T_12976; // @[LoadQueue.scala 141:18:@11780.4]
  wire  entriesToCheck_5_7; // @[LoadQueue.scala 141:26:@11781.4]
  wire  _T_12978; // @[LoadQueue.scala 141:18:@11782.4]
  wire  entriesToCheck_5_8; // @[LoadQueue.scala 141:26:@11783.4]
  wire  _T_12980; // @[LoadQueue.scala 141:18:@11784.4]
  wire  entriesToCheck_5_9; // @[LoadQueue.scala 141:26:@11785.4]
  wire  _T_12982; // @[LoadQueue.scala 141:18:@11786.4]
  wire  entriesToCheck_5_10; // @[LoadQueue.scala 141:26:@11787.4]
  wire  _T_12984; // @[LoadQueue.scala 141:18:@11788.4]
  wire  entriesToCheck_5_11; // @[LoadQueue.scala 141:26:@11789.4]
  wire  _T_12986; // @[LoadQueue.scala 141:18:@11790.4]
  wire  entriesToCheck_5_12; // @[LoadQueue.scala 141:26:@11791.4]
  wire  _T_12988; // @[LoadQueue.scala 141:18:@11792.4]
  wire  entriesToCheck_5_13; // @[LoadQueue.scala 141:26:@11793.4]
  wire  _T_12990; // @[LoadQueue.scala 141:18:@11794.4]
  wire  entriesToCheck_5_14; // @[LoadQueue.scala 141:26:@11795.4]
  wire  _T_12992; // @[LoadQueue.scala 141:18:@11796.4]
  wire  entriesToCheck_5_15; // @[LoadQueue.scala 141:26:@11797.4]
  wire  _T_12994; // @[LoadQueue.scala 141:18:@11814.4]
  wire  entriesToCheck_6_0; // @[LoadQueue.scala 141:26:@11815.4]
  wire  _T_12996; // @[LoadQueue.scala 141:18:@11816.4]
  wire  entriesToCheck_6_1; // @[LoadQueue.scala 141:26:@11817.4]
  wire  _T_12998; // @[LoadQueue.scala 141:18:@11818.4]
  wire  entriesToCheck_6_2; // @[LoadQueue.scala 141:26:@11819.4]
  wire  _T_13000; // @[LoadQueue.scala 141:18:@11820.4]
  wire  entriesToCheck_6_3; // @[LoadQueue.scala 141:26:@11821.4]
  wire  _T_13002; // @[LoadQueue.scala 141:18:@11822.4]
  wire  entriesToCheck_6_4; // @[LoadQueue.scala 141:26:@11823.4]
  wire  _T_13004; // @[LoadQueue.scala 141:18:@11824.4]
  wire  entriesToCheck_6_5; // @[LoadQueue.scala 141:26:@11825.4]
  wire  _T_13006; // @[LoadQueue.scala 141:18:@11826.4]
  wire  entriesToCheck_6_6; // @[LoadQueue.scala 141:26:@11827.4]
  wire  _T_13008; // @[LoadQueue.scala 141:18:@11828.4]
  wire  entriesToCheck_6_7; // @[LoadQueue.scala 141:26:@11829.4]
  wire  _T_13010; // @[LoadQueue.scala 141:18:@11830.4]
  wire  entriesToCheck_6_8; // @[LoadQueue.scala 141:26:@11831.4]
  wire  _T_13012; // @[LoadQueue.scala 141:18:@11832.4]
  wire  entriesToCheck_6_9; // @[LoadQueue.scala 141:26:@11833.4]
  wire  _T_13014; // @[LoadQueue.scala 141:18:@11834.4]
  wire  entriesToCheck_6_10; // @[LoadQueue.scala 141:26:@11835.4]
  wire  _T_13016; // @[LoadQueue.scala 141:18:@11836.4]
  wire  entriesToCheck_6_11; // @[LoadQueue.scala 141:26:@11837.4]
  wire  _T_13018; // @[LoadQueue.scala 141:18:@11838.4]
  wire  entriesToCheck_6_12; // @[LoadQueue.scala 141:26:@11839.4]
  wire  _T_13020; // @[LoadQueue.scala 141:18:@11840.4]
  wire  entriesToCheck_6_13; // @[LoadQueue.scala 141:26:@11841.4]
  wire  _T_13022; // @[LoadQueue.scala 141:18:@11842.4]
  wire  entriesToCheck_6_14; // @[LoadQueue.scala 141:26:@11843.4]
  wire  _T_13024; // @[LoadQueue.scala 141:18:@11844.4]
  wire  entriesToCheck_6_15; // @[LoadQueue.scala 141:26:@11845.4]
  wire  _T_13026; // @[LoadQueue.scala 141:18:@11862.4]
  wire  entriesToCheck_7_0; // @[LoadQueue.scala 141:26:@11863.4]
  wire  _T_13028; // @[LoadQueue.scala 141:18:@11864.4]
  wire  entriesToCheck_7_1; // @[LoadQueue.scala 141:26:@11865.4]
  wire  _T_13030; // @[LoadQueue.scala 141:18:@11866.4]
  wire  entriesToCheck_7_2; // @[LoadQueue.scala 141:26:@11867.4]
  wire  _T_13032; // @[LoadQueue.scala 141:18:@11868.4]
  wire  entriesToCheck_7_3; // @[LoadQueue.scala 141:26:@11869.4]
  wire  _T_13034; // @[LoadQueue.scala 141:18:@11870.4]
  wire  entriesToCheck_7_4; // @[LoadQueue.scala 141:26:@11871.4]
  wire  _T_13036; // @[LoadQueue.scala 141:18:@11872.4]
  wire  entriesToCheck_7_5; // @[LoadQueue.scala 141:26:@11873.4]
  wire  _T_13038; // @[LoadQueue.scala 141:18:@11874.4]
  wire  entriesToCheck_7_6; // @[LoadQueue.scala 141:26:@11875.4]
  wire  _T_13040; // @[LoadQueue.scala 141:18:@11876.4]
  wire  entriesToCheck_7_7; // @[LoadQueue.scala 141:26:@11877.4]
  wire  _T_13042; // @[LoadQueue.scala 141:18:@11878.4]
  wire  entriesToCheck_7_8; // @[LoadQueue.scala 141:26:@11879.4]
  wire  _T_13044; // @[LoadQueue.scala 141:18:@11880.4]
  wire  entriesToCheck_7_9; // @[LoadQueue.scala 141:26:@11881.4]
  wire  _T_13046; // @[LoadQueue.scala 141:18:@11882.4]
  wire  entriesToCheck_7_10; // @[LoadQueue.scala 141:26:@11883.4]
  wire  _T_13048; // @[LoadQueue.scala 141:18:@11884.4]
  wire  entriesToCheck_7_11; // @[LoadQueue.scala 141:26:@11885.4]
  wire  _T_13050; // @[LoadQueue.scala 141:18:@11886.4]
  wire  entriesToCheck_7_12; // @[LoadQueue.scala 141:26:@11887.4]
  wire  _T_13052; // @[LoadQueue.scala 141:18:@11888.4]
  wire  entriesToCheck_7_13; // @[LoadQueue.scala 141:26:@11889.4]
  wire  _T_13054; // @[LoadQueue.scala 141:18:@11890.4]
  wire  entriesToCheck_7_14; // @[LoadQueue.scala 141:26:@11891.4]
  wire  _T_13056; // @[LoadQueue.scala 141:18:@11892.4]
  wire  entriesToCheck_7_15; // @[LoadQueue.scala 141:26:@11893.4]
  wire  _T_13058; // @[LoadQueue.scala 141:18:@11910.4]
  wire  entriesToCheck_8_0; // @[LoadQueue.scala 141:26:@11911.4]
  wire  _T_13060; // @[LoadQueue.scala 141:18:@11912.4]
  wire  entriesToCheck_8_1; // @[LoadQueue.scala 141:26:@11913.4]
  wire  _T_13062; // @[LoadQueue.scala 141:18:@11914.4]
  wire  entriesToCheck_8_2; // @[LoadQueue.scala 141:26:@11915.4]
  wire  _T_13064; // @[LoadQueue.scala 141:18:@11916.4]
  wire  entriesToCheck_8_3; // @[LoadQueue.scala 141:26:@11917.4]
  wire  _T_13066; // @[LoadQueue.scala 141:18:@11918.4]
  wire  entriesToCheck_8_4; // @[LoadQueue.scala 141:26:@11919.4]
  wire  _T_13068; // @[LoadQueue.scala 141:18:@11920.4]
  wire  entriesToCheck_8_5; // @[LoadQueue.scala 141:26:@11921.4]
  wire  _T_13070; // @[LoadQueue.scala 141:18:@11922.4]
  wire  entriesToCheck_8_6; // @[LoadQueue.scala 141:26:@11923.4]
  wire  _T_13072; // @[LoadQueue.scala 141:18:@11924.4]
  wire  entriesToCheck_8_7; // @[LoadQueue.scala 141:26:@11925.4]
  wire  _T_13074; // @[LoadQueue.scala 141:18:@11926.4]
  wire  entriesToCheck_8_8; // @[LoadQueue.scala 141:26:@11927.4]
  wire  _T_13076; // @[LoadQueue.scala 141:18:@11928.4]
  wire  entriesToCheck_8_9; // @[LoadQueue.scala 141:26:@11929.4]
  wire  _T_13078; // @[LoadQueue.scala 141:18:@11930.4]
  wire  entriesToCheck_8_10; // @[LoadQueue.scala 141:26:@11931.4]
  wire  _T_13080; // @[LoadQueue.scala 141:18:@11932.4]
  wire  entriesToCheck_8_11; // @[LoadQueue.scala 141:26:@11933.4]
  wire  _T_13082; // @[LoadQueue.scala 141:18:@11934.4]
  wire  entriesToCheck_8_12; // @[LoadQueue.scala 141:26:@11935.4]
  wire  _T_13084; // @[LoadQueue.scala 141:18:@11936.4]
  wire  entriesToCheck_8_13; // @[LoadQueue.scala 141:26:@11937.4]
  wire  _T_13086; // @[LoadQueue.scala 141:18:@11938.4]
  wire  entriesToCheck_8_14; // @[LoadQueue.scala 141:26:@11939.4]
  wire  _T_13088; // @[LoadQueue.scala 141:18:@11940.4]
  wire  entriesToCheck_8_15; // @[LoadQueue.scala 141:26:@11941.4]
  wire  _T_13090; // @[LoadQueue.scala 141:18:@11958.4]
  wire  entriesToCheck_9_0; // @[LoadQueue.scala 141:26:@11959.4]
  wire  _T_13092; // @[LoadQueue.scala 141:18:@11960.4]
  wire  entriesToCheck_9_1; // @[LoadQueue.scala 141:26:@11961.4]
  wire  _T_13094; // @[LoadQueue.scala 141:18:@11962.4]
  wire  entriesToCheck_9_2; // @[LoadQueue.scala 141:26:@11963.4]
  wire  _T_13096; // @[LoadQueue.scala 141:18:@11964.4]
  wire  entriesToCheck_9_3; // @[LoadQueue.scala 141:26:@11965.4]
  wire  _T_13098; // @[LoadQueue.scala 141:18:@11966.4]
  wire  entriesToCheck_9_4; // @[LoadQueue.scala 141:26:@11967.4]
  wire  _T_13100; // @[LoadQueue.scala 141:18:@11968.4]
  wire  entriesToCheck_9_5; // @[LoadQueue.scala 141:26:@11969.4]
  wire  _T_13102; // @[LoadQueue.scala 141:18:@11970.4]
  wire  entriesToCheck_9_6; // @[LoadQueue.scala 141:26:@11971.4]
  wire  _T_13104; // @[LoadQueue.scala 141:18:@11972.4]
  wire  entriesToCheck_9_7; // @[LoadQueue.scala 141:26:@11973.4]
  wire  _T_13106; // @[LoadQueue.scala 141:18:@11974.4]
  wire  entriesToCheck_9_8; // @[LoadQueue.scala 141:26:@11975.4]
  wire  _T_13108; // @[LoadQueue.scala 141:18:@11976.4]
  wire  entriesToCheck_9_9; // @[LoadQueue.scala 141:26:@11977.4]
  wire  _T_13110; // @[LoadQueue.scala 141:18:@11978.4]
  wire  entriesToCheck_9_10; // @[LoadQueue.scala 141:26:@11979.4]
  wire  _T_13112; // @[LoadQueue.scala 141:18:@11980.4]
  wire  entriesToCheck_9_11; // @[LoadQueue.scala 141:26:@11981.4]
  wire  _T_13114; // @[LoadQueue.scala 141:18:@11982.4]
  wire  entriesToCheck_9_12; // @[LoadQueue.scala 141:26:@11983.4]
  wire  _T_13116; // @[LoadQueue.scala 141:18:@11984.4]
  wire  entriesToCheck_9_13; // @[LoadQueue.scala 141:26:@11985.4]
  wire  _T_13118; // @[LoadQueue.scala 141:18:@11986.4]
  wire  entriesToCheck_9_14; // @[LoadQueue.scala 141:26:@11987.4]
  wire  _T_13120; // @[LoadQueue.scala 141:18:@11988.4]
  wire  entriesToCheck_9_15; // @[LoadQueue.scala 141:26:@11989.4]
  wire  _T_13122; // @[LoadQueue.scala 141:18:@12006.4]
  wire  entriesToCheck_10_0; // @[LoadQueue.scala 141:26:@12007.4]
  wire  _T_13124; // @[LoadQueue.scala 141:18:@12008.4]
  wire  entriesToCheck_10_1; // @[LoadQueue.scala 141:26:@12009.4]
  wire  _T_13126; // @[LoadQueue.scala 141:18:@12010.4]
  wire  entriesToCheck_10_2; // @[LoadQueue.scala 141:26:@12011.4]
  wire  _T_13128; // @[LoadQueue.scala 141:18:@12012.4]
  wire  entriesToCheck_10_3; // @[LoadQueue.scala 141:26:@12013.4]
  wire  _T_13130; // @[LoadQueue.scala 141:18:@12014.4]
  wire  entriesToCheck_10_4; // @[LoadQueue.scala 141:26:@12015.4]
  wire  _T_13132; // @[LoadQueue.scala 141:18:@12016.4]
  wire  entriesToCheck_10_5; // @[LoadQueue.scala 141:26:@12017.4]
  wire  _T_13134; // @[LoadQueue.scala 141:18:@12018.4]
  wire  entriesToCheck_10_6; // @[LoadQueue.scala 141:26:@12019.4]
  wire  _T_13136; // @[LoadQueue.scala 141:18:@12020.4]
  wire  entriesToCheck_10_7; // @[LoadQueue.scala 141:26:@12021.4]
  wire  _T_13138; // @[LoadQueue.scala 141:18:@12022.4]
  wire  entriesToCheck_10_8; // @[LoadQueue.scala 141:26:@12023.4]
  wire  _T_13140; // @[LoadQueue.scala 141:18:@12024.4]
  wire  entriesToCheck_10_9; // @[LoadQueue.scala 141:26:@12025.4]
  wire  _T_13142; // @[LoadQueue.scala 141:18:@12026.4]
  wire  entriesToCheck_10_10; // @[LoadQueue.scala 141:26:@12027.4]
  wire  _T_13144; // @[LoadQueue.scala 141:18:@12028.4]
  wire  entriesToCheck_10_11; // @[LoadQueue.scala 141:26:@12029.4]
  wire  _T_13146; // @[LoadQueue.scala 141:18:@12030.4]
  wire  entriesToCheck_10_12; // @[LoadQueue.scala 141:26:@12031.4]
  wire  _T_13148; // @[LoadQueue.scala 141:18:@12032.4]
  wire  entriesToCheck_10_13; // @[LoadQueue.scala 141:26:@12033.4]
  wire  _T_13150; // @[LoadQueue.scala 141:18:@12034.4]
  wire  entriesToCheck_10_14; // @[LoadQueue.scala 141:26:@12035.4]
  wire  _T_13152; // @[LoadQueue.scala 141:18:@12036.4]
  wire  entriesToCheck_10_15; // @[LoadQueue.scala 141:26:@12037.4]
  wire  _T_13154; // @[LoadQueue.scala 141:18:@12054.4]
  wire  entriesToCheck_11_0; // @[LoadQueue.scala 141:26:@12055.4]
  wire  _T_13156; // @[LoadQueue.scala 141:18:@12056.4]
  wire  entriesToCheck_11_1; // @[LoadQueue.scala 141:26:@12057.4]
  wire  _T_13158; // @[LoadQueue.scala 141:18:@12058.4]
  wire  entriesToCheck_11_2; // @[LoadQueue.scala 141:26:@12059.4]
  wire  _T_13160; // @[LoadQueue.scala 141:18:@12060.4]
  wire  entriesToCheck_11_3; // @[LoadQueue.scala 141:26:@12061.4]
  wire  _T_13162; // @[LoadQueue.scala 141:18:@12062.4]
  wire  entriesToCheck_11_4; // @[LoadQueue.scala 141:26:@12063.4]
  wire  _T_13164; // @[LoadQueue.scala 141:18:@12064.4]
  wire  entriesToCheck_11_5; // @[LoadQueue.scala 141:26:@12065.4]
  wire  _T_13166; // @[LoadQueue.scala 141:18:@12066.4]
  wire  entriesToCheck_11_6; // @[LoadQueue.scala 141:26:@12067.4]
  wire  _T_13168; // @[LoadQueue.scala 141:18:@12068.4]
  wire  entriesToCheck_11_7; // @[LoadQueue.scala 141:26:@12069.4]
  wire  _T_13170; // @[LoadQueue.scala 141:18:@12070.4]
  wire  entriesToCheck_11_8; // @[LoadQueue.scala 141:26:@12071.4]
  wire  _T_13172; // @[LoadQueue.scala 141:18:@12072.4]
  wire  entriesToCheck_11_9; // @[LoadQueue.scala 141:26:@12073.4]
  wire  _T_13174; // @[LoadQueue.scala 141:18:@12074.4]
  wire  entriesToCheck_11_10; // @[LoadQueue.scala 141:26:@12075.4]
  wire  _T_13176; // @[LoadQueue.scala 141:18:@12076.4]
  wire  entriesToCheck_11_11; // @[LoadQueue.scala 141:26:@12077.4]
  wire  _T_13178; // @[LoadQueue.scala 141:18:@12078.4]
  wire  entriesToCheck_11_12; // @[LoadQueue.scala 141:26:@12079.4]
  wire  _T_13180; // @[LoadQueue.scala 141:18:@12080.4]
  wire  entriesToCheck_11_13; // @[LoadQueue.scala 141:26:@12081.4]
  wire  _T_13182; // @[LoadQueue.scala 141:18:@12082.4]
  wire  entriesToCheck_11_14; // @[LoadQueue.scala 141:26:@12083.4]
  wire  _T_13184; // @[LoadQueue.scala 141:18:@12084.4]
  wire  entriesToCheck_11_15; // @[LoadQueue.scala 141:26:@12085.4]
  wire  _T_13186; // @[LoadQueue.scala 141:18:@12102.4]
  wire  entriesToCheck_12_0; // @[LoadQueue.scala 141:26:@12103.4]
  wire  _T_13188; // @[LoadQueue.scala 141:18:@12104.4]
  wire  entriesToCheck_12_1; // @[LoadQueue.scala 141:26:@12105.4]
  wire  _T_13190; // @[LoadQueue.scala 141:18:@12106.4]
  wire  entriesToCheck_12_2; // @[LoadQueue.scala 141:26:@12107.4]
  wire  _T_13192; // @[LoadQueue.scala 141:18:@12108.4]
  wire  entriesToCheck_12_3; // @[LoadQueue.scala 141:26:@12109.4]
  wire  _T_13194; // @[LoadQueue.scala 141:18:@12110.4]
  wire  entriesToCheck_12_4; // @[LoadQueue.scala 141:26:@12111.4]
  wire  _T_13196; // @[LoadQueue.scala 141:18:@12112.4]
  wire  entriesToCheck_12_5; // @[LoadQueue.scala 141:26:@12113.4]
  wire  _T_13198; // @[LoadQueue.scala 141:18:@12114.4]
  wire  entriesToCheck_12_6; // @[LoadQueue.scala 141:26:@12115.4]
  wire  _T_13200; // @[LoadQueue.scala 141:18:@12116.4]
  wire  entriesToCheck_12_7; // @[LoadQueue.scala 141:26:@12117.4]
  wire  _T_13202; // @[LoadQueue.scala 141:18:@12118.4]
  wire  entriesToCheck_12_8; // @[LoadQueue.scala 141:26:@12119.4]
  wire  _T_13204; // @[LoadQueue.scala 141:18:@12120.4]
  wire  entriesToCheck_12_9; // @[LoadQueue.scala 141:26:@12121.4]
  wire  _T_13206; // @[LoadQueue.scala 141:18:@12122.4]
  wire  entriesToCheck_12_10; // @[LoadQueue.scala 141:26:@12123.4]
  wire  _T_13208; // @[LoadQueue.scala 141:18:@12124.4]
  wire  entriesToCheck_12_11; // @[LoadQueue.scala 141:26:@12125.4]
  wire  _T_13210; // @[LoadQueue.scala 141:18:@12126.4]
  wire  entriesToCheck_12_12; // @[LoadQueue.scala 141:26:@12127.4]
  wire  _T_13212; // @[LoadQueue.scala 141:18:@12128.4]
  wire  entriesToCheck_12_13; // @[LoadQueue.scala 141:26:@12129.4]
  wire  _T_13214; // @[LoadQueue.scala 141:18:@12130.4]
  wire  entriesToCheck_12_14; // @[LoadQueue.scala 141:26:@12131.4]
  wire  _T_13216; // @[LoadQueue.scala 141:18:@12132.4]
  wire  entriesToCheck_12_15; // @[LoadQueue.scala 141:26:@12133.4]
  wire  _T_13218; // @[LoadQueue.scala 141:18:@12150.4]
  wire  entriesToCheck_13_0; // @[LoadQueue.scala 141:26:@12151.4]
  wire  _T_13220; // @[LoadQueue.scala 141:18:@12152.4]
  wire  entriesToCheck_13_1; // @[LoadQueue.scala 141:26:@12153.4]
  wire  _T_13222; // @[LoadQueue.scala 141:18:@12154.4]
  wire  entriesToCheck_13_2; // @[LoadQueue.scala 141:26:@12155.4]
  wire  _T_13224; // @[LoadQueue.scala 141:18:@12156.4]
  wire  entriesToCheck_13_3; // @[LoadQueue.scala 141:26:@12157.4]
  wire  _T_13226; // @[LoadQueue.scala 141:18:@12158.4]
  wire  entriesToCheck_13_4; // @[LoadQueue.scala 141:26:@12159.4]
  wire  _T_13228; // @[LoadQueue.scala 141:18:@12160.4]
  wire  entriesToCheck_13_5; // @[LoadQueue.scala 141:26:@12161.4]
  wire  _T_13230; // @[LoadQueue.scala 141:18:@12162.4]
  wire  entriesToCheck_13_6; // @[LoadQueue.scala 141:26:@12163.4]
  wire  _T_13232; // @[LoadQueue.scala 141:18:@12164.4]
  wire  entriesToCheck_13_7; // @[LoadQueue.scala 141:26:@12165.4]
  wire  _T_13234; // @[LoadQueue.scala 141:18:@12166.4]
  wire  entriesToCheck_13_8; // @[LoadQueue.scala 141:26:@12167.4]
  wire  _T_13236; // @[LoadQueue.scala 141:18:@12168.4]
  wire  entriesToCheck_13_9; // @[LoadQueue.scala 141:26:@12169.4]
  wire  _T_13238; // @[LoadQueue.scala 141:18:@12170.4]
  wire  entriesToCheck_13_10; // @[LoadQueue.scala 141:26:@12171.4]
  wire  _T_13240; // @[LoadQueue.scala 141:18:@12172.4]
  wire  entriesToCheck_13_11; // @[LoadQueue.scala 141:26:@12173.4]
  wire  _T_13242; // @[LoadQueue.scala 141:18:@12174.4]
  wire  entriesToCheck_13_12; // @[LoadQueue.scala 141:26:@12175.4]
  wire  _T_13244; // @[LoadQueue.scala 141:18:@12176.4]
  wire  entriesToCheck_13_13; // @[LoadQueue.scala 141:26:@12177.4]
  wire  _T_13246; // @[LoadQueue.scala 141:18:@12178.4]
  wire  entriesToCheck_13_14; // @[LoadQueue.scala 141:26:@12179.4]
  wire  _T_13248; // @[LoadQueue.scala 141:18:@12180.4]
  wire  entriesToCheck_13_15; // @[LoadQueue.scala 141:26:@12181.4]
  wire  _T_13250; // @[LoadQueue.scala 141:18:@12198.4]
  wire  entriesToCheck_14_0; // @[LoadQueue.scala 141:26:@12199.4]
  wire  _T_13252; // @[LoadQueue.scala 141:18:@12200.4]
  wire  entriesToCheck_14_1; // @[LoadQueue.scala 141:26:@12201.4]
  wire  _T_13254; // @[LoadQueue.scala 141:18:@12202.4]
  wire  entriesToCheck_14_2; // @[LoadQueue.scala 141:26:@12203.4]
  wire  _T_13256; // @[LoadQueue.scala 141:18:@12204.4]
  wire  entriesToCheck_14_3; // @[LoadQueue.scala 141:26:@12205.4]
  wire  _T_13258; // @[LoadQueue.scala 141:18:@12206.4]
  wire  entriesToCheck_14_4; // @[LoadQueue.scala 141:26:@12207.4]
  wire  _T_13260; // @[LoadQueue.scala 141:18:@12208.4]
  wire  entriesToCheck_14_5; // @[LoadQueue.scala 141:26:@12209.4]
  wire  _T_13262; // @[LoadQueue.scala 141:18:@12210.4]
  wire  entriesToCheck_14_6; // @[LoadQueue.scala 141:26:@12211.4]
  wire  _T_13264; // @[LoadQueue.scala 141:18:@12212.4]
  wire  entriesToCheck_14_7; // @[LoadQueue.scala 141:26:@12213.4]
  wire  _T_13266; // @[LoadQueue.scala 141:18:@12214.4]
  wire  entriesToCheck_14_8; // @[LoadQueue.scala 141:26:@12215.4]
  wire  _T_13268; // @[LoadQueue.scala 141:18:@12216.4]
  wire  entriesToCheck_14_9; // @[LoadQueue.scala 141:26:@12217.4]
  wire  _T_13270; // @[LoadQueue.scala 141:18:@12218.4]
  wire  entriesToCheck_14_10; // @[LoadQueue.scala 141:26:@12219.4]
  wire  _T_13272; // @[LoadQueue.scala 141:18:@12220.4]
  wire  entriesToCheck_14_11; // @[LoadQueue.scala 141:26:@12221.4]
  wire  _T_13274; // @[LoadQueue.scala 141:18:@12222.4]
  wire  entriesToCheck_14_12; // @[LoadQueue.scala 141:26:@12223.4]
  wire  _T_13276; // @[LoadQueue.scala 141:18:@12224.4]
  wire  entriesToCheck_14_13; // @[LoadQueue.scala 141:26:@12225.4]
  wire  _T_13278; // @[LoadQueue.scala 141:18:@12226.4]
  wire  entriesToCheck_14_14; // @[LoadQueue.scala 141:26:@12227.4]
  wire  _T_13280; // @[LoadQueue.scala 141:18:@12228.4]
  wire  entriesToCheck_14_15; // @[LoadQueue.scala 141:26:@12229.4]
  wire  _T_13282; // @[LoadQueue.scala 141:18:@12246.4]
  wire  entriesToCheck_15_0; // @[LoadQueue.scala 141:26:@12247.4]
  wire  _T_13284; // @[LoadQueue.scala 141:18:@12248.4]
  wire  entriesToCheck_15_1; // @[LoadQueue.scala 141:26:@12249.4]
  wire  _T_13286; // @[LoadQueue.scala 141:18:@12250.4]
  wire  entriesToCheck_15_2; // @[LoadQueue.scala 141:26:@12251.4]
  wire  _T_13288; // @[LoadQueue.scala 141:18:@12252.4]
  wire  entriesToCheck_15_3; // @[LoadQueue.scala 141:26:@12253.4]
  wire  _T_13290; // @[LoadQueue.scala 141:18:@12254.4]
  wire  entriesToCheck_15_4; // @[LoadQueue.scala 141:26:@12255.4]
  wire  _T_13292; // @[LoadQueue.scala 141:18:@12256.4]
  wire  entriesToCheck_15_5; // @[LoadQueue.scala 141:26:@12257.4]
  wire  _T_13294; // @[LoadQueue.scala 141:18:@12258.4]
  wire  entriesToCheck_15_6; // @[LoadQueue.scala 141:26:@12259.4]
  wire  _T_13296; // @[LoadQueue.scala 141:18:@12260.4]
  wire  entriesToCheck_15_7; // @[LoadQueue.scala 141:26:@12261.4]
  wire  _T_13298; // @[LoadQueue.scala 141:18:@12262.4]
  wire  entriesToCheck_15_8; // @[LoadQueue.scala 141:26:@12263.4]
  wire  _T_13300; // @[LoadQueue.scala 141:18:@12264.4]
  wire  entriesToCheck_15_9; // @[LoadQueue.scala 141:26:@12265.4]
  wire  _T_13302; // @[LoadQueue.scala 141:18:@12266.4]
  wire  entriesToCheck_15_10; // @[LoadQueue.scala 141:26:@12267.4]
  wire  _T_13304; // @[LoadQueue.scala 141:18:@12268.4]
  wire  entriesToCheck_15_11; // @[LoadQueue.scala 141:26:@12269.4]
  wire  _T_13306; // @[LoadQueue.scala 141:18:@12270.4]
  wire  entriesToCheck_15_12; // @[LoadQueue.scala 141:26:@12271.4]
  wire  _T_13308; // @[LoadQueue.scala 141:18:@12272.4]
  wire  entriesToCheck_15_13; // @[LoadQueue.scala 141:26:@12273.4]
  wire  _T_13310; // @[LoadQueue.scala 141:18:@12274.4]
  wire  entriesToCheck_15_14; // @[LoadQueue.scala 141:26:@12275.4]
  wire  _T_13312; // @[LoadQueue.scala 141:18:@12276.4]
  wire  entriesToCheck_15_15; // @[LoadQueue.scala 141:26:@12277.4]
  wire  _T_14544; // @[LoadQueue.scala 151:92:@12295.4]
  wire  _T_14545; // @[LoadQueue.scala 152:41:@12296.4]
  wire  _T_14546; // @[LoadQueue.scala 153:30:@12297.4]
  wire  conflict_0_0; // @[LoadQueue.scala 152:68:@12298.4]
  wire  _T_14548; // @[LoadQueue.scala 151:92:@12300.4]
  wire  _T_14549; // @[LoadQueue.scala 152:41:@12301.4]
  wire  _T_14550; // @[LoadQueue.scala 153:30:@12302.4]
  wire  conflict_0_1; // @[LoadQueue.scala 152:68:@12303.4]
  wire  _T_14552; // @[LoadQueue.scala 151:92:@12305.4]
  wire  _T_14553; // @[LoadQueue.scala 152:41:@12306.4]
  wire  _T_14554; // @[LoadQueue.scala 153:30:@12307.4]
  wire  conflict_0_2; // @[LoadQueue.scala 152:68:@12308.4]
  wire  _T_14556; // @[LoadQueue.scala 151:92:@12310.4]
  wire  _T_14557; // @[LoadQueue.scala 152:41:@12311.4]
  wire  _T_14558; // @[LoadQueue.scala 153:30:@12312.4]
  wire  conflict_0_3; // @[LoadQueue.scala 152:68:@12313.4]
  wire  _T_14560; // @[LoadQueue.scala 151:92:@12315.4]
  wire  _T_14561; // @[LoadQueue.scala 152:41:@12316.4]
  wire  _T_14562; // @[LoadQueue.scala 153:30:@12317.4]
  wire  conflict_0_4; // @[LoadQueue.scala 152:68:@12318.4]
  wire  _T_14564; // @[LoadQueue.scala 151:92:@12320.4]
  wire  _T_14565; // @[LoadQueue.scala 152:41:@12321.4]
  wire  _T_14566; // @[LoadQueue.scala 153:30:@12322.4]
  wire  conflict_0_5; // @[LoadQueue.scala 152:68:@12323.4]
  wire  _T_14568; // @[LoadQueue.scala 151:92:@12325.4]
  wire  _T_14569; // @[LoadQueue.scala 152:41:@12326.4]
  wire  _T_14570; // @[LoadQueue.scala 153:30:@12327.4]
  wire  conflict_0_6; // @[LoadQueue.scala 152:68:@12328.4]
  wire  _T_14572; // @[LoadQueue.scala 151:92:@12330.4]
  wire  _T_14573; // @[LoadQueue.scala 152:41:@12331.4]
  wire  _T_14574; // @[LoadQueue.scala 153:30:@12332.4]
  wire  conflict_0_7; // @[LoadQueue.scala 152:68:@12333.4]
  wire  _T_14576; // @[LoadQueue.scala 151:92:@12335.4]
  wire  _T_14577; // @[LoadQueue.scala 152:41:@12336.4]
  wire  _T_14578; // @[LoadQueue.scala 153:30:@12337.4]
  wire  conflict_0_8; // @[LoadQueue.scala 152:68:@12338.4]
  wire  _T_14580; // @[LoadQueue.scala 151:92:@12340.4]
  wire  _T_14581; // @[LoadQueue.scala 152:41:@12341.4]
  wire  _T_14582; // @[LoadQueue.scala 153:30:@12342.4]
  wire  conflict_0_9; // @[LoadQueue.scala 152:68:@12343.4]
  wire  _T_14584; // @[LoadQueue.scala 151:92:@12345.4]
  wire  _T_14585; // @[LoadQueue.scala 152:41:@12346.4]
  wire  _T_14586; // @[LoadQueue.scala 153:30:@12347.4]
  wire  conflict_0_10; // @[LoadQueue.scala 152:68:@12348.4]
  wire  _T_14588; // @[LoadQueue.scala 151:92:@12350.4]
  wire  _T_14589; // @[LoadQueue.scala 152:41:@12351.4]
  wire  _T_14590; // @[LoadQueue.scala 153:30:@12352.4]
  wire  conflict_0_11; // @[LoadQueue.scala 152:68:@12353.4]
  wire  _T_14592; // @[LoadQueue.scala 151:92:@12355.4]
  wire  _T_14593; // @[LoadQueue.scala 152:41:@12356.4]
  wire  _T_14594; // @[LoadQueue.scala 153:30:@12357.4]
  wire  conflict_0_12; // @[LoadQueue.scala 152:68:@12358.4]
  wire  _T_14596; // @[LoadQueue.scala 151:92:@12360.4]
  wire  _T_14597; // @[LoadQueue.scala 152:41:@12361.4]
  wire  _T_14598; // @[LoadQueue.scala 153:30:@12362.4]
  wire  conflict_0_13; // @[LoadQueue.scala 152:68:@12363.4]
  wire  _T_14600; // @[LoadQueue.scala 151:92:@12365.4]
  wire  _T_14601; // @[LoadQueue.scala 152:41:@12366.4]
  wire  _T_14602; // @[LoadQueue.scala 153:30:@12367.4]
  wire  conflict_0_14; // @[LoadQueue.scala 152:68:@12368.4]
  wire  _T_14604; // @[LoadQueue.scala 151:92:@12370.4]
  wire  _T_14605; // @[LoadQueue.scala 152:41:@12371.4]
  wire  _T_14606; // @[LoadQueue.scala 153:30:@12372.4]
  wire  conflict_0_15; // @[LoadQueue.scala 152:68:@12373.4]
  wire  _T_14608; // @[LoadQueue.scala 151:92:@12375.4]
  wire  _T_14609; // @[LoadQueue.scala 152:41:@12376.4]
  wire  _T_14610; // @[LoadQueue.scala 153:30:@12377.4]
  wire  conflict_1_0; // @[LoadQueue.scala 152:68:@12378.4]
  wire  _T_14612; // @[LoadQueue.scala 151:92:@12380.4]
  wire  _T_14613; // @[LoadQueue.scala 152:41:@12381.4]
  wire  _T_14614; // @[LoadQueue.scala 153:30:@12382.4]
  wire  conflict_1_1; // @[LoadQueue.scala 152:68:@12383.4]
  wire  _T_14616; // @[LoadQueue.scala 151:92:@12385.4]
  wire  _T_14617; // @[LoadQueue.scala 152:41:@12386.4]
  wire  _T_14618; // @[LoadQueue.scala 153:30:@12387.4]
  wire  conflict_1_2; // @[LoadQueue.scala 152:68:@12388.4]
  wire  _T_14620; // @[LoadQueue.scala 151:92:@12390.4]
  wire  _T_14621; // @[LoadQueue.scala 152:41:@12391.4]
  wire  _T_14622; // @[LoadQueue.scala 153:30:@12392.4]
  wire  conflict_1_3; // @[LoadQueue.scala 152:68:@12393.4]
  wire  _T_14624; // @[LoadQueue.scala 151:92:@12395.4]
  wire  _T_14625; // @[LoadQueue.scala 152:41:@12396.4]
  wire  _T_14626; // @[LoadQueue.scala 153:30:@12397.4]
  wire  conflict_1_4; // @[LoadQueue.scala 152:68:@12398.4]
  wire  _T_14628; // @[LoadQueue.scala 151:92:@12400.4]
  wire  _T_14629; // @[LoadQueue.scala 152:41:@12401.4]
  wire  _T_14630; // @[LoadQueue.scala 153:30:@12402.4]
  wire  conflict_1_5; // @[LoadQueue.scala 152:68:@12403.4]
  wire  _T_14632; // @[LoadQueue.scala 151:92:@12405.4]
  wire  _T_14633; // @[LoadQueue.scala 152:41:@12406.4]
  wire  _T_14634; // @[LoadQueue.scala 153:30:@12407.4]
  wire  conflict_1_6; // @[LoadQueue.scala 152:68:@12408.4]
  wire  _T_14636; // @[LoadQueue.scala 151:92:@12410.4]
  wire  _T_14637; // @[LoadQueue.scala 152:41:@12411.4]
  wire  _T_14638; // @[LoadQueue.scala 153:30:@12412.4]
  wire  conflict_1_7; // @[LoadQueue.scala 152:68:@12413.4]
  wire  _T_14640; // @[LoadQueue.scala 151:92:@12415.4]
  wire  _T_14641; // @[LoadQueue.scala 152:41:@12416.4]
  wire  _T_14642; // @[LoadQueue.scala 153:30:@12417.4]
  wire  conflict_1_8; // @[LoadQueue.scala 152:68:@12418.4]
  wire  _T_14644; // @[LoadQueue.scala 151:92:@12420.4]
  wire  _T_14645; // @[LoadQueue.scala 152:41:@12421.4]
  wire  _T_14646; // @[LoadQueue.scala 153:30:@12422.4]
  wire  conflict_1_9; // @[LoadQueue.scala 152:68:@12423.4]
  wire  _T_14648; // @[LoadQueue.scala 151:92:@12425.4]
  wire  _T_14649; // @[LoadQueue.scala 152:41:@12426.4]
  wire  _T_14650; // @[LoadQueue.scala 153:30:@12427.4]
  wire  conflict_1_10; // @[LoadQueue.scala 152:68:@12428.4]
  wire  _T_14652; // @[LoadQueue.scala 151:92:@12430.4]
  wire  _T_14653; // @[LoadQueue.scala 152:41:@12431.4]
  wire  _T_14654; // @[LoadQueue.scala 153:30:@12432.4]
  wire  conflict_1_11; // @[LoadQueue.scala 152:68:@12433.4]
  wire  _T_14656; // @[LoadQueue.scala 151:92:@12435.4]
  wire  _T_14657; // @[LoadQueue.scala 152:41:@12436.4]
  wire  _T_14658; // @[LoadQueue.scala 153:30:@12437.4]
  wire  conflict_1_12; // @[LoadQueue.scala 152:68:@12438.4]
  wire  _T_14660; // @[LoadQueue.scala 151:92:@12440.4]
  wire  _T_14661; // @[LoadQueue.scala 152:41:@12441.4]
  wire  _T_14662; // @[LoadQueue.scala 153:30:@12442.4]
  wire  conflict_1_13; // @[LoadQueue.scala 152:68:@12443.4]
  wire  _T_14664; // @[LoadQueue.scala 151:92:@12445.4]
  wire  _T_14665; // @[LoadQueue.scala 152:41:@12446.4]
  wire  _T_14666; // @[LoadQueue.scala 153:30:@12447.4]
  wire  conflict_1_14; // @[LoadQueue.scala 152:68:@12448.4]
  wire  _T_14668; // @[LoadQueue.scala 151:92:@12450.4]
  wire  _T_14669; // @[LoadQueue.scala 152:41:@12451.4]
  wire  _T_14670; // @[LoadQueue.scala 153:30:@12452.4]
  wire  conflict_1_15; // @[LoadQueue.scala 152:68:@12453.4]
  wire  _T_14672; // @[LoadQueue.scala 151:92:@12455.4]
  wire  _T_14673; // @[LoadQueue.scala 152:41:@12456.4]
  wire  _T_14674; // @[LoadQueue.scala 153:30:@12457.4]
  wire  conflict_2_0; // @[LoadQueue.scala 152:68:@12458.4]
  wire  _T_14676; // @[LoadQueue.scala 151:92:@12460.4]
  wire  _T_14677; // @[LoadQueue.scala 152:41:@12461.4]
  wire  _T_14678; // @[LoadQueue.scala 153:30:@12462.4]
  wire  conflict_2_1; // @[LoadQueue.scala 152:68:@12463.4]
  wire  _T_14680; // @[LoadQueue.scala 151:92:@12465.4]
  wire  _T_14681; // @[LoadQueue.scala 152:41:@12466.4]
  wire  _T_14682; // @[LoadQueue.scala 153:30:@12467.4]
  wire  conflict_2_2; // @[LoadQueue.scala 152:68:@12468.4]
  wire  _T_14684; // @[LoadQueue.scala 151:92:@12470.4]
  wire  _T_14685; // @[LoadQueue.scala 152:41:@12471.4]
  wire  _T_14686; // @[LoadQueue.scala 153:30:@12472.4]
  wire  conflict_2_3; // @[LoadQueue.scala 152:68:@12473.4]
  wire  _T_14688; // @[LoadQueue.scala 151:92:@12475.4]
  wire  _T_14689; // @[LoadQueue.scala 152:41:@12476.4]
  wire  _T_14690; // @[LoadQueue.scala 153:30:@12477.4]
  wire  conflict_2_4; // @[LoadQueue.scala 152:68:@12478.4]
  wire  _T_14692; // @[LoadQueue.scala 151:92:@12480.4]
  wire  _T_14693; // @[LoadQueue.scala 152:41:@12481.4]
  wire  _T_14694; // @[LoadQueue.scala 153:30:@12482.4]
  wire  conflict_2_5; // @[LoadQueue.scala 152:68:@12483.4]
  wire  _T_14696; // @[LoadQueue.scala 151:92:@12485.4]
  wire  _T_14697; // @[LoadQueue.scala 152:41:@12486.4]
  wire  _T_14698; // @[LoadQueue.scala 153:30:@12487.4]
  wire  conflict_2_6; // @[LoadQueue.scala 152:68:@12488.4]
  wire  _T_14700; // @[LoadQueue.scala 151:92:@12490.4]
  wire  _T_14701; // @[LoadQueue.scala 152:41:@12491.4]
  wire  _T_14702; // @[LoadQueue.scala 153:30:@12492.4]
  wire  conflict_2_7; // @[LoadQueue.scala 152:68:@12493.4]
  wire  _T_14704; // @[LoadQueue.scala 151:92:@12495.4]
  wire  _T_14705; // @[LoadQueue.scala 152:41:@12496.4]
  wire  _T_14706; // @[LoadQueue.scala 153:30:@12497.4]
  wire  conflict_2_8; // @[LoadQueue.scala 152:68:@12498.4]
  wire  _T_14708; // @[LoadQueue.scala 151:92:@12500.4]
  wire  _T_14709; // @[LoadQueue.scala 152:41:@12501.4]
  wire  _T_14710; // @[LoadQueue.scala 153:30:@12502.4]
  wire  conflict_2_9; // @[LoadQueue.scala 152:68:@12503.4]
  wire  _T_14712; // @[LoadQueue.scala 151:92:@12505.4]
  wire  _T_14713; // @[LoadQueue.scala 152:41:@12506.4]
  wire  _T_14714; // @[LoadQueue.scala 153:30:@12507.4]
  wire  conflict_2_10; // @[LoadQueue.scala 152:68:@12508.4]
  wire  _T_14716; // @[LoadQueue.scala 151:92:@12510.4]
  wire  _T_14717; // @[LoadQueue.scala 152:41:@12511.4]
  wire  _T_14718; // @[LoadQueue.scala 153:30:@12512.4]
  wire  conflict_2_11; // @[LoadQueue.scala 152:68:@12513.4]
  wire  _T_14720; // @[LoadQueue.scala 151:92:@12515.4]
  wire  _T_14721; // @[LoadQueue.scala 152:41:@12516.4]
  wire  _T_14722; // @[LoadQueue.scala 153:30:@12517.4]
  wire  conflict_2_12; // @[LoadQueue.scala 152:68:@12518.4]
  wire  _T_14724; // @[LoadQueue.scala 151:92:@12520.4]
  wire  _T_14725; // @[LoadQueue.scala 152:41:@12521.4]
  wire  _T_14726; // @[LoadQueue.scala 153:30:@12522.4]
  wire  conflict_2_13; // @[LoadQueue.scala 152:68:@12523.4]
  wire  _T_14728; // @[LoadQueue.scala 151:92:@12525.4]
  wire  _T_14729; // @[LoadQueue.scala 152:41:@12526.4]
  wire  _T_14730; // @[LoadQueue.scala 153:30:@12527.4]
  wire  conflict_2_14; // @[LoadQueue.scala 152:68:@12528.4]
  wire  _T_14732; // @[LoadQueue.scala 151:92:@12530.4]
  wire  _T_14733; // @[LoadQueue.scala 152:41:@12531.4]
  wire  _T_14734; // @[LoadQueue.scala 153:30:@12532.4]
  wire  conflict_2_15; // @[LoadQueue.scala 152:68:@12533.4]
  wire  _T_14736; // @[LoadQueue.scala 151:92:@12535.4]
  wire  _T_14737; // @[LoadQueue.scala 152:41:@12536.4]
  wire  _T_14738; // @[LoadQueue.scala 153:30:@12537.4]
  wire  conflict_3_0; // @[LoadQueue.scala 152:68:@12538.4]
  wire  _T_14740; // @[LoadQueue.scala 151:92:@12540.4]
  wire  _T_14741; // @[LoadQueue.scala 152:41:@12541.4]
  wire  _T_14742; // @[LoadQueue.scala 153:30:@12542.4]
  wire  conflict_3_1; // @[LoadQueue.scala 152:68:@12543.4]
  wire  _T_14744; // @[LoadQueue.scala 151:92:@12545.4]
  wire  _T_14745; // @[LoadQueue.scala 152:41:@12546.4]
  wire  _T_14746; // @[LoadQueue.scala 153:30:@12547.4]
  wire  conflict_3_2; // @[LoadQueue.scala 152:68:@12548.4]
  wire  _T_14748; // @[LoadQueue.scala 151:92:@12550.4]
  wire  _T_14749; // @[LoadQueue.scala 152:41:@12551.4]
  wire  _T_14750; // @[LoadQueue.scala 153:30:@12552.4]
  wire  conflict_3_3; // @[LoadQueue.scala 152:68:@12553.4]
  wire  _T_14752; // @[LoadQueue.scala 151:92:@12555.4]
  wire  _T_14753; // @[LoadQueue.scala 152:41:@12556.4]
  wire  _T_14754; // @[LoadQueue.scala 153:30:@12557.4]
  wire  conflict_3_4; // @[LoadQueue.scala 152:68:@12558.4]
  wire  _T_14756; // @[LoadQueue.scala 151:92:@12560.4]
  wire  _T_14757; // @[LoadQueue.scala 152:41:@12561.4]
  wire  _T_14758; // @[LoadQueue.scala 153:30:@12562.4]
  wire  conflict_3_5; // @[LoadQueue.scala 152:68:@12563.4]
  wire  _T_14760; // @[LoadQueue.scala 151:92:@12565.4]
  wire  _T_14761; // @[LoadQueue.scala 152:41:@12566.4]
  wire  _T_14762; // @[LoadQueue.scala 153:30:@12567.4]
  wire  conflict_3_6; // @[LoadQueue.scala 152:68:@12568.4]
  wire  _T_14764; // @[LoadQueue.scala 151:92:@12570.4]
  wire  _T_14765; // @[LoadQueue.scala 152:41:@12571.4]
  wire  _T_14766; // @[LoadQueue.scala 153:30:@12572.4]
  wire  conflict_3_7; // @[LoadQueue.scala 152:68:@12573.4]
  wire  _T_14768; // @[LoadQueue.scala 151:92:@12575.4]
  wire  _T_14769; // @[LoadQueue.scala 152:41:@12576.4]
  wire  _T_14770; // @[LoadQueue.scala 153:30:@12577.4]
  wire  conflict_3_8; // @[LoadQueue.scala 152:68:@12578.4]
  wire  _T_14772; // @[LoadQueue.scala 151:92:@12580.4]
  wire  _T_14773; // @[LoadQueue.scala 152:41:@12581.4]
  wire  _T_14774; // @[LoadQueue.scala 153:30:@12582.4]
  wire  conflict_3_9; // @[LoadQueue.scala 152:68:@12583.4]
  wire  _T_14776; // @[LoadQueue.scala 151:92:@12585.4]
  wire  _T_14777; // @[LoadQueue.scala 152:41:@12586.4]
  wire  _T_14778; // @[LoadQueue.scala 153:30:@12587.4]
  wire  conflict_3_10; // @[LoadQueue.scala 152:68:@12588.4]
  wire  _T_14780; // @[LoadQueue.scala 151:92:@12590.4]
  wire  _T_14781; // @[LoadQueue.scala 152:41:@12591.4]
  wire  _T_14782; // @[LoadQueue.scala 153:30:@12592.4]
  wire  conflict_3_11; // @[LoadQueue.scala 152:68:@12593.4]
  wire  _T_14784; // @[LoadQueue.scala 151:92:@12595.4]
  wire  _T_14785; // @[LoadQueue.scala 152:41:@12596.4]
  wire  _T_14786; // @[LoadQueue.scala 153:30:@12597.4]
  wire  conflict_3_12; // @[LoadQueue.scala 152:68:@12598.4]
  wire  _T_14788; // @[LoadQueue.scala 151:92:@12600.4]
  wire  _T_14789; // @[LoadQueue.scala 152:41:@12601.4]
  wire  _T_14790; // @[LoadQueue.scala 153:30:@12602.4]
  wire  conflict_3_13; // @[LoadQueue.scala 152:68:@12603.4]
  wire  _T_14792; // @[LoadQueue.scala 151:92:@12605.4]
  wire  _T_14793; // @[LoadQueue.scala 152:41:@12606.4]
  wire  _T_14794; // @[LoadQueue.scala 153:30:@12607.4]
  wire  conflict_3_14; // @[LoadQueue.scala 152:68:@12608.4]
  wire  _T_14796; // @[LoadQueue.scala 151:92:@12610.4]
  wire  _T_14797; // @[LoadQueue.scala 152:41:@12611.4]
  wire  _T_14798; // @[LoadQueue.scala 153:30:@12612.4]
  wire  conflict_3_15; // @[LoadQueue.scala 152:68:@12613.4]
  wire  _T_14800; // @[LoadQueue.scala 151:92:@12615.4]
  wire  _T_14801; // @[LoadQueue.scala 152:41:@12616.4]
  wire  _T_14802; // @[LoadQueue.scala 153:30:@12617.4]
  wire  conflict_4_0; // @[LoadQueue.scala 152:68:@12618.4]
  wire  _T_14804; // @[LoadQueue.scala 151:92:@12620.4]
  wire  _T_14805; // @[LoadQueue.scala 152:41:@12621.4]
  wire  _T_14806; // @[LoadQueue.scala 153:30:@12622.4]
  wire  conflict_4_1; // @[LoadQueue.scala 152:68:@12623.4]
  wire  _T_14808; // @[LoadQueue.scala 151:92:@12625.4]
  wire  _T_14809; // @[LoadQueue.scala 152:41:@12626.4]
  wire  _T_14810; // @[LoadQueue.scala 153:30:@12627.4]
  wire  conflict_4_2; // @[LoadQueue.scala 152:68:@12628.4]
  wire  _T_14812; // @[LoadQueue.scala 151:92:@12630.4]
  wire  _T_14813; // @[LoadQueue.scala 152:41:@12631.4]
  wire  _T_14814; // @[LoadQueue.scala 153:30:@12632.4]
  wire  conflict_4_3; // @[LoadQueue.scala 152:68:@12633.4]
  wire  _T_14816; // @[LoadQueue.scala 151:92:@12635.4]
  wire  _T_14817; // @[LoadQueue.scala 152:41:@12636.4]
  wire  _T_14818; // @[LoadQueue.scala 153:30:@12637.4]
  wire  conflict_4_4; // @[LoadQueue.scala 152:68:@12638.4]
  wire  _T_14820; // @[LoadQueue.scala 151:92:@12640.4]
  wire  _T_14821; // @[LoadQueue.scala 152:41:@12641.4]
  wire  _T_14822; // @[LoadQueue.scala 153:30:@12642.4]
  wire  conflict_4_5; // @[LoadQueue.scala 152:68:@12643.4]
  wire  _T_14824; // @[LoadQueue.scala 151:92:@12645.4]
  wire  _T_14825; // @[LoadQueue.scala 152:41:@12646.4]
  wire  _T_14826; // @[LoadQueue.scala 153:30:@12647.4]
  wire  conflict_4_6; // @[LoadQueue.scala 152:68:@12648.4]
  wire  _T_14828; // @[LoadQueue.scala 151:92:@12650.4]
  wire  _T_14829; // @[LoadQueue.scala 152:41:@12651.4]
  wire  _T_14830; // @[LoadQueue.scala 153:30:@12652.4]
  wire  conflict_4_7; // @[LoadQueue.scala 152:68:@12653.4]
  wire  _T_14832; // @[LoadQueue.scala 151:92:@12655.4]
  wire  _T_14833; // @[LoadQueue.scala 152:41:@12656.4]
  wire  _T_14834; // @[LoadQueue.scala 153:30:@12657.4]
  wire  conflict_4_8; // @[LoadQueue.scala 152:68:@12658.4]
  wire  _T_14836; // @[LoadQueue.scala 151:92:@12660.4]
  wire  _T_14837; // @[LoadQueue.scala 152:41:@12661.4]
  wire  _T_14838; // @[LoadQueue.scala 153:30:@12662.4]
  wire  conflict_4_9; // @[LoadQueue.scala 152:68:@12663.4]
  wire  _T_14840; // @[LoadQueue.scala 151:92:@12665.4]
  wire  _T_14841; // @[LoadQueue.scala 152:41:@12666.4]
  wire  _T_14842; // @[LoadQueue.scala 153:30:@12667.4]
  wire  conflict_4_10; // @[LoadQueue.scala 152:68:@12668.4]
  wire  _T_14844; // @[LoadQueue.scala 151:92:@12670.4]
  wire  _T_14845; // @[LoadQueue.scala 152:41:@12671.4]
  wire  _T_14846; // @[LoadQueue.scala 153:30:@12672.4]
  wire  conflict_4_11; // @[LoadQueue.scala 152:68:@12673.4]
  wire  _T_14848; // @[LoadQueue.scala 151:92:@12675.4]
  wire  _T_14849; // @[LoadQueue.scala 152:41:@12676.4]
  wire  _T_14850; // @[LoadQueue.scala 153:30:@12677.4]
  wire  conflict_4_12; // @[LoadQueue.scala 152:68:@12678.4]
  wire  _T_14852; // @[LoadQueue.scala 151:92:@12680.4]
  wire  _T_14853; // @[LoadQueue.scala 152:41:@12681.4]
  wire  _T_14854; // @[LoadQueue.scala 153:30:@12682.4]
  wire  conflict_4_13; // @[LoadQueue.scala 152:68:@12683.4]
  wire  _T_14856; // @[LoadQueue.scala 151:92:@12685.4]
  wire  _T_14857; // @[LoadQueue.scala 152:41:@12686.4]
  wire  _T_14858; // @[LoadQueue.scala 153:30:@12687.4]
  wire  conflict_4_14; // @[LoadQueue.scala 152:68:@12688.4]
  wire  _T_14860; // @[LoadQueue.scala 151:92:@12690.4]
  wire  _T_14861; // @[LoadQueue.scala 152:41:@12691.4]
  wire  _T_14862; // @[LoadQueue.scala 153:30:@12692.4]
  wire  conflict_4_15; // @[LoadQueue.scala 152:68:@12693.4]
  wire  _T_14864; // @[LoadQueue.scala 151:92:@12695.4]
  wire  _T_14865; // @[LoadQueue.scala 152:41:@12696.4]
  wire  _T_14866; // @[LoadQueue.scala 153:30:@12697.4]
  wire  conflict_5_0; // @[LoadQueue.scala 152:68:@12698.4]
  wire  _T_14868; // @[LoadQueue.scala 151:92:@12700.4]
  wire  _T_14869; // @[LoadQueue.scala 152:41:@12701.4]
  wire  _T_14870; // @[LoadQueue.scala 153:30:@12702.4]
  wire  conflict_5_1; // @[LoadQueue.scala 152:68:@12703.4]
  wire  _T_14872; // @[LoadQueue.scala 151:92:@12705.4]
  wire  _T_14873; // @[LoadQueue.scala 152:41:@12706.4]
  wire  _T_14874; // @[LoadQueue.scala 153:30:@12707.4]
  wire  conflict_5_2; // @[LoadQueue.scala 152:68:@12708.4]
  wire  _T_14876; // @[LoadQueue.scala 151:92:@12710.4]
  wire  _T_14877; // @[LoadQueue.scala 152:41:@12711.4]
  wire  _T_14878; // @[LoadQueue.scala 153:30:@12712.4]
  wire  conflict_5_3; // @[LoadQueue.scala 152:68:@12713.4]
  wire  _T_14880; // @[LoadQueue.scala 151:92:@12715.4]
  wire  _T_14881; // @[LoadQueue.scala 152:41:@12716.4]
  wire  _T_14882; // @[LoadQueue.scala 153:30:@12717.4]
  wire  conflict_5_4; // @[LoadQueue.scala 152:68:@12718.4]
  wire  _T_14884; // @[LoadQueue.scala 151:92:@12720.4]
  wire  _T_14885; // @[LoadQueue.scala 152:41:@12721.4]
  wire  _T_14886; // @[LoadQueue.scala 153:30:@12722.4]
  wire  conflict_5_5; // @[LoadQueue.scala 152:68:@12723.4]
  wire  _T_14888; // @[LoadQueue.scala 151:92:@12725.4]
  wire  _T_14889; // @[LoadQueue.scala 152:41:@12726.4]
  wire  _T_14890; // @[LoadQueue.scala 153:30:@12727.4]
  wire  conflict_5_6; // @[LoadQueue.scala 152:68:@12728.4]
  wire  _T_14892; // @[LoadQueue.scala 151:92:@12730.4]
  wire  _T_14893; // @[LoadQueue.scala 152:41:@12731.4]
  wire  _T_14894; // @[LoadQueue.scala 153:30:@12732.4]
  wire  conflict_5_7; // @[LoadQueue.scala 152:68:@12733.4]
  wire  _T_14896; // @[LoadQueue.scala 151:92:@12735.4]
  wire  _T_14897; // @[LoadQueue.scala 152:41:@12736.4]
  wire  _T_14898; // @[LoadQueue.scala 153:30:@12737.4]
  wire  conflict_5_8; // @[LoadQueue.scala 152:68:@12738.4]
  wire  _T_14900; // @[LoadQueue.scala 151:92:@12740.4]
  wire  _T_14901; // @[LoadQueue.scala 152:41:@12741.4]
  wire  _T_14902; // @[LoadQueue.scala 153:30:@12742.4]
  wire  conflict_5_9; // @[LoadQueue.scala 152:68:@12743.4]
  wire  _T_14904; // @[LoadQueue.scala 151:92:@12745.4]
  wire  _T_14905; // @[LoadQueue.scala 152:41:@12746.4]
  wire  _T_14906; // @[LoadQueue.scala 153:30:@12747.4]
  wire  conflict_5_10; // @[LoadQueue.scala 152:68:@12748.4]
  wire  _T_14908; // @[LoadQueue.scala 151:92:@12750.4]
  wire  _T_14909; // @[LoadQueue.scala 152:41:@12751.4]
  wire  _T_14910; // @[LoadQueue.scala 153:30:@12752.4]
  wire  conflict_5_11; // @[LoadQueue.scala 152:68:@12753.4]
  wire  _T_14912; // @[LoadQueue.scala 151:92:@12755.4]
  wire  _T_14913; // @[LoadQueue.scala 152:41:@12756.4]
  wire  _T_14914; // @[LoadQueue.scala 153:30:@12757.4]
  wire  conflict_5_12; // @[LoadQueue.scala 152:68:@12758.4]
  wire  _T_14916; // @[LoadQueue.scala 151:92:@12760.4]
  wire  _T_14917; // @[LoadQueue.scala 152:41:@12761.4]
  wire  _T_14918; // @[LoadQueue.scala 153:30:@12762.4]
  wire  conflict_5_13; // @[LoadQueue.scala 152:68:@12763.4]
  wire  _T_14920; // @[LoadQueue.scala 151:92:@12765.4]
  wire  _T_14921; // @[LoadQueue.scala 152:41:@12766.4]
  wire  _T_14922; // @[LoadQueue.scala 153:30:@12767.4]
  wire  conflict_5_14; // @[LoadQueue.scala 152:68:@12768.4]
  wire  _T_14924; // @[LoadQueue.scala 151:92:@12770.4]
  wire  _T_14925; // @[LoadQueue.scala 152:41:@12771.4]
  wire  _T_14926; // @[LoadQueue.scala 153:30:@12772.4]
  wire  conflict_5_15; // @[LoadQueue.scala 152:68:@12773.4]
  wire  _T_14928; // @[LoadQueue.scala 151:92:@12775.4]
  wire  _T_14929; // @[LoadQueue.scala 152:41:@12776.4]
  wire  _T_14930; // @[LoadQueue.scala 153:30:@12777.4]
  wire  conflict_6_0; // @[LoadQueue.scala 152:68:@12778.4]
  wire  _T_14932; // @[LoadQueue.scala 151:92:@12780.4]
  wire  _T_14933; // @[LoadQueue.scala 152:41:@12781.4]
  wire  _T_14934; // @[LoadQueue.scala 153:30:@12782.4]
  wire  conflict_6_1; // @[LoadQueue.scala 152:68:@12783.4]
  wire  _T_14936; // @[LoadQueue.scala 151:92:@12785.4]
  wire  _T_14937; // @[LoadQueue.scala 152:41:@12786.4]
  wire  _T_14938; // @[LoadQueue.scala 153:30:@12787.4]
  wire  conflict_6_2; // @[LoadQueue.scala 152:68:@12788.4]
  wire  _T_14940; // @[LoadQueue.scala 151:92:@12790.4]
  wire  _T_14941; // @[LoadQueue.scala 152:41:@12791.4]
  wire  _T_14942; // @[LoadQueue.scala 153:30:@12792.4]
  wire  conflict_6_3; // @[LoadQueue.scala 152:68:@12793.4]
  wire  _T_14944; // @[LoadQueue.scala 151:92:@12795.4]
  wire  _T_14945; // @[LoadQueue.scala 152:41:@12796.4]
  wire  _T_14946; // @[LoadQueue.scala 153:30:@12797.4]
  wire  conflict_6_4; // @[LoadQueue.scala 152:68:@12798.4]
  wire  _T_14948; // @[LoadQueue.scala 151:92:@12800.4]
  wire  _T_14949; // @[LoadQueue.scala 152:41:@12801.4]
  wire  _T_14950; // @[LoadQueue.scala 153:30:@12802.4]
  wire  conflict_6_5; // @[LoadQueue.scala 152:68:@12803.4]
  wire  _T_14952; // @[LoadQueue.scala 151:92:@12805.4]
  wire  _T_14953; // @[LoadQueue.scala 152:41:@12806.4]
  wire  _T_14954; // @[LoadQueue.scala 153:30:@12807.4]
  wire  conflict_6_6; // @[LoadQueue.scala 152:68:@12808.4]
  wire  _T_14956; // @[LoadQueue.scala 151:92:@12810.4]
  wire  _T_14957; // @[LoadQueue.scala 152:41:@12811.4]
  wire  _T_14958; // @[LoadQueue.scala 153:30:@12812.4]
  wire  conflict_6_7; // @[LoadQueue.scala 152:68:@12813.4]
  wire  _T_14960; // @[LoadQueue.scala 151:92:@12815.4]
  wire  _T_14961; // @[LoadQueue.scala 152:41:@12816.4]
  wire  _T_14962; // @[LoadQueue.scala 153:30:@12817.4]
  wire  conflict_6_8; // @[LoadQueue.scala 152:68:@12818.4]
  wire  _T_14964; // @[LoadQueue.scala 151:92:@12820.4]
  wire  _T_14965; // @[LoadQueue.scala 152:41:@12821.4]
  wire  _T_14966; // @[LoadQueue.scala 153:30:@12822.4]
  wire  conflict_6_9; // @[LoadQueue.scala 152:68:@12823.4]
  wire  _T_14968; // @[LoadQueue.scala 151:92:@12825.4]
  wire  _T_14969; // @[LoadQueue.scala 152:41:@12826.4]
  wire  _T_14970; // @[LoadQueue.scala 153:30:@12827.4]
  wire  conflict_6_10; // @[LoadQueue.scala 152:68:@12828.4]
  wire  _T_14972; // @[LoadQueue.scala 151:92:@12830.4]
  wire  _T_14973; // @[LoadQueue.scala 152:41:@12831.4]
  wire  _T_14974; // @[LoadQueue.scala 153:30:@12832.4]
  wire  conflict_6_11; // @[LoadQueue.scala 152:68:@12833.4]
  wire  _T_14976; // @[LoadQueue.scala 151:92:@12835.4]
  wire  _T_14977; // @[LoadQueue.scala 152:41:@12836.4]
  wire  _T_14978; // @[LoadQueue.scala 153:30:@12837.4]
  wire  conflict_6_12; // @[LoadQueue.scala 152:68:@12838.4]
  wire  _T_14980; // @[LoadQueue.scala 151:92:@12840.4]
  wire  _T_14981; // @[LoadQueue.scala 152:41:@12841.4]
  wire  _T_14982; // @[LoadQueue.scala 153:30:@12842.4]
  wire  conflict_6_13; // @[LoadQueue.scala 152:68:@12843.4]
  wire  _T_14984; // @[LoadQueue.scala 151:92:@12845.4]
  wire  _T_14985; // @[LoadQueue.scala 152:41:@12846.4]
  wire  _T_14986; // @[LoadQueue.scala 153:30:@12847.4]
  wire  conflict_6_14; // @[LoadQueue.scala 152:68:@12848.4]
  wire  _T_14988; // @[LoadQueue.scala 151:92:@12850.4]
  wire  _T_14989; // @[LoadQueue.scala 152:41:@12851.4]
  wire  _T_14990; // @[LoadQueue.scala 153:30:@12852.4]
  wire  conflict_6_15; // @[LoadQueue.scala 152:68:@12853.4]
  wire  _T_14992; // @[LoadQueue.scala 151:92:@12855.4]
  wire  _T_14993; // @[LoadQueue.scala 152:41:@12856.4]
  wire  _T_14994; // @[LoadQueue.scala 153:30:@12857.4]
  wire  conflict_7_0; // @[LoadQueue.scala 152:68:@12858.4]
  wire  _T_14996; // @[LoadQueue.scala 151:92:@12860.4]
  wire  _T_14997; // @[LoadQueue.scala 152:41:@12861.4]
  wire  _T_14998; // @[LoadQueue.scala 153:30:@12862.4]
  wire  conflict_7_1; // @[LoadQueue.scala 152:68:@12863.4]
  wire  _T_15000; // @[LoadQueue.scala 151:92:@12865.4]
  wire  _T_15001; // @[LoadQueue.scala 152:41:@12866.4]
  wire  _T_15002; // @[LoadQueue.scala 153:30:@12867.4]
  wire  conflict_7_2; // @[LoadQueue.scala 152:68:@12868.4]
  wire  _T_15004; // @[LoadQueue.scala 151:92:@12870.4]
  wire  _T_15005; // @[LoadQueue.scala 152:41:@12871.4]
  wire  _T_15006; // @[LoadQueue.scala 153:30:@12872.4]
  wire  conflict_7_3; // @[LoadQueue.scala 152:68:@12873.4]
  wire  _T_15008; // @[LoadQueue.scala 151:92:@12875.4]
  wire  _T_15009; // @[LoadQueue.scala 152:41:@12876.4]
  wire  _T_15010; // @[LoadQueue.scala 153:30:@12877.4]
  wire  conflict_7_4; // @[LoadQueue.scala 152:68:@12878.4]
  wire  _T_15012; // @[LoadQueue.scala 151:92:@12880.4]
  wire  _T_15013; // @[LoadQueue.scala 152:41:@12881.4]
  wire  _T_15014; // @[LoadQueue.scala 153:30:@12882.4]
  wire  conflict_7_5; // @[LoadQueue.scala 152:68:@12883.4]
  wire  _T_15016; // @[LoadQueue.scala 151:92:@12885.4]
  wire  _T_15017; // @[LoadQueue.scala 152:41:@12886.4]
  wire  _T_15018; // @[LoadQueue.scala 153:30:@12887.4]
  wire  conflict_7_6; // @[LoadQueue.scala 152:68:@12888.4]
  wire  _T_15020; // @[LoadQueue.scala 151:92:@12890.4]
  wire  _T_15021; // @[LoadQueue.scala 152:41:@12891.4]
  wire  _T_15022; // @[LoadQueue.scala 153:30:@12892.4]
  wire  conflict_7_7; // @[LoadQueue.scala 152:68:@12893.4]
  wire  _T_15024; // @[LoadQueue.scala 151:92:@12895.4]
  wire  _T_15025; // @[LoadQueue.scala 152:41:@12896.4]
  wire  _T_15026; // @[LoadQueue.scala 153:30:@12897.4]
  wire  conflict_7_8; // @[LoadQueue.scala 152:68:@12898.4]
  wire  _T_15028; // @[LoadQueue.scala 151:92:@12900.4]
  wire  _T_15029; // @[LoadQueue.scala 152:41:@12901.4]
  wire  _T_15030; // @[LoadQueue.scala 153:30:@12902.4]
  wire  conflict_7_9; // @[LoadQueue.scala 152:68:@12903.4]
  wire  _T_15032; // @[LoadQueue.scala 151:92:@12905.4]
  wire  _T_15033; // @[LoadQueue.scala 152:41:@12906.4]
  wire  _T_15034; // @[LoadQueue.scala 153:30:@12907.4]
  wire  conflict_7_10; // @[LoadQueue.scala 152:68:@12908.4]
  wire  _T_15036; // @[LoadQueue.scala 151:92:@12910.4]
  wire  _T_15037; // @[LoadQueue.scala 152:41:@12911.4]
  wire  _T_15038; // @[LoadQueue.scala 153:30:@12912.4]
  wire  conflict_7_11; // @[LoadQueue.scala 152:68:@12913.4]
  wire  _T_15040; // @[LoadQueue.scala 151:92:@12915.4]
  wire  _T_15041; // @[LoadQueue.scala 152:41:@12916.4]
  wire  _T_15042; // @[LoadQueue.scala 153:30:@12917.4]
  wire  conflict_7_12; // @[LoadQueue.scala 152:68:@12918.4]
  wire  _T_15044; // @[LoadQueue.scala 151:92:@12920.4]
  wire  _T_15045; // @[LoadQueue.scala 152:41:@12921.4]
  wire  _T_15046; // @[LoadQueue.scala 153:30:@12922.4]
  wire  conflict_7_13; // @[LoadQueue.scala 152:68:@12923.4]
  wire  _T_15048; // @[LoadQueue.scala 151:92:@12925.4]
  wire  _T_15049; // @[LoadQueue.scala 152:41:@12926.4]
  wire  _T_15050; // @[LoadQueue.scala 153:30:@12927.4]
  wire  conflict_7_14; // @[LoadQueue.scala 152:68:@12928.4]
  wire  _T_15052; // @[LoadQueue.scala 151:92:@12930.4]
  wire  _T_15053; // @[LoadQueue.scala 152:41:@12931.4]
  wire  _T_15054; // @[LoadQueue.scala 153:30:@12932.4]
  wire  conflict_7_15; // @[LoadQueue.scala 152:68:@12933.4]
  wire  _T_15056; // @[LoadQueue.scala 151:92:@12935.4]
  wire  _T_15057; // @[LoadQueue.scala 152:41:@12936.4]
  wire  _T_15058; // @[LoadQueue.scala 153:30:@12937.4]
  wire  conflict_8_0; // @[LoadQueue.scala 152:68:@12938.4]
  wire  _T_15060; // @[LoadQueue.scala 151:92:@12940.4]
  wire  _T_15061; // @[LoadQueue.scala 152:41:@12941.4]
  wire  _T_15062; // @[LoadQueue.scala 153:30:@12942.4]
  wire  conflict_8_1; // @[LoadQueue.scala 152:68:@12943.4]
  wire  _T_15064; // @[LoadQueue.scala 151:92:@12945.4]
  wire  _T_15065; // @[LoadQueue.scala 152:41:@12946.4]
  wire  _T_15066; // @[LoadQueue.scala 153:30:@12947.4]
  wire  conflict_8_2; // @[LoadQueue.scala 152:68:@12948.4]
  wire  _T_15068; // @[LoadQueue.scala 151:92:@12950.4]
  wire  _T_15069; // @[LoadQueue.scala 152:41:@12951.4]
  wire  _T_15070; // @[LoadQueue.scala 153:30:@12952.4]
  wire  conflict_8_3; // @[LoadQueue.scala 152:68:@12953.4]
  wire  _T_15072; // @[LoadQueue.scala 151:92:@12955.4]
  wire  _T_15073; // @[LoadQueue.scala 152:41:@12956.4]
  wire  _T_15074; // @[LoadQueue.scala 153:30:@12957.4]
  wire  conflict_8_4; // @[LoadQueue.scala 152:68:@12958.4]
  wire  _T_15076; // @[LoadQueue.scala 151:92:@12960.4]
  wire  _T_15077; // @[LoadQueue.scala 152:41:@12961.4]
  wire  _T_15078; // @[LoadQueue.scala 153:30:@12962.4]
  wire  conflict_8_5; // @[LoadQueue.scala 152:68:@12963.4]
  wire  _T_15080; // @[LoadQueue.scala 151:92:@12965.4]
  wire  _T_15081; // @[LoadQueue.scala 152:41:@12966.4]
  wire  _T_15082; // @[LoadQueue.scala 153:30:@12967.4]
  wire  conflict_8_6; // @[LoadQueue.scala 152:68:@12968.4]
  wire  _T_15084; // @[LoadQueue.scala 151:92:@12970.4]
  wire  _T_15085; // @[LoadQueue.scala 152:41:@12971.4]
  wire  _T_15086; // @[LoadQueue.scala 153:30:@12972.4]
  wire  conflict_8_7; // @[LoadQueue.scala 152:68:@12973.4]
  wire  _T_15088; // @[LoadQueue.scala 151:92:@12975.4]
  wire  _T_15089; // @[LoadQueue.scala 152:41:@12976.4]
  wire  _T_15090; // @[LoadQueue.scala 153:30:@12977.4]
  wire  conflict_8_8; // @[LoadQueue.scala 152:68:@12978.4]
  wire  _T_15092; // @[LoadQueue.scala 151:92:@12980.4]
  wire  _T_15093; // @[LoadQueue.scala 152:41:@12981.4]
  wire  _T_15094; // @[LoadQueue.scala 153:30:@12982.4]
  wire  conflict_8_9; // @[LoadQueue.scala 152:68:@12983.4]
  wire  _T_15096; // @[LoadQueue.scala 151:92:@12985.4]
  wire  _T_15097; // @[LoadQueue.scala 152:41:@12986.4]
  wire  _T_15098; // @[LoadQueue.scala 153:30:@12987.4]
  wire  conflict_8_10; // @[LoadQueue.scala 152:68:@12988.4]
  wire  _T_15100; // @[LoadQueue.scala 151:92:@12990.4]
  wire  _T_15101; // @[LoadQueue.scala 152:41:@12991.4]
  wire  _T_15102; // @[LoadQueue.scala 153:30:@12992.4]
  wire  conflict_8_11; // @[LoadQueue.scala 152:68:@12993.4]
  wire  _T_15104; // @[LoadQueue.scala 151:92:@12995.4]
  wire  _T_15105; // @[LoadQueue.scala 152:41:@12996.4]
  wire  _T_15106; // @[LoadQueue.scala 153:30:@12997.4]
  wire  conflict_8_12; // @[LoadQueue.scala 152:68:@12998.4]
  wire  _T_15108; // @[LoadQueue.scala 151:92:@13000.4]
  wire  _T_15109; // @[LoadQueue.scala 152:41:@13001.4]
  wire  _T_15110; // @[LoadQueue.scala 153:30:@13002.4]
  wire  conflict_8_13; // @[LoadQueue.scala 152:68:@13003.4]
  wire  _T_15112; // @[LoadQueue.scala 151:92:@13005.4]
  wire  _T_15113; // @[LoadQueue.scala 152:41:@13006.4]
  wire  _T_15114; // @[LoadQueue.scala 153:30:@13007.4]
  wire  conflict_8_14; // @[LoadQueue.scala 152:68:@13008.4]
  wire  _T_15116; // @[LoadQueue.scala 151:92:@13010.4]
  wire  _T_15117; // @[LoadQueue.scala 152:41:@13011.4]
  wire  _T_15118; // @[LoadQueue.scala 153:30:@13012.4]
  wire  conflict_8_15; // @[LoadQueue.scala 152:68:@13013.4]
  wire  _T_15120; // @[LoadQueue.scala 151:92:@13015.4]
  wire  _T_15121; // @[LoadQueue.scala 152:41:@13016.4]
  wire  _T_15122; // @[LoadQueue.scala 153:30:@13017.4]
  wire  conflict_9_0; // @[LoadQueue.scala 152:68:@13018.4]
  wire  _T_15124; // @[LoadQueue.scala 151:92:@13020.4]
  wire  _T_15125; // @[LoadQueue.scala 152:41:@13021.4]
  wire  _T_15126; // @[LoadQueue.scala 153:30:@13022.4]
  wire  conflict_9_1; // @[LoadQueue.scala 152:68:@13023.4]
  wire  _T_15128; // @[LoadQueue.scala 151:92:@13025.4]
  wire  _T_15129; // @[LoadQueue.scala 152:41:@13026.4]
  wire  _T_15130; // @[LoadQueue.scala 153:30:@13027.4]
  wire  conflict_9_2; // @[LoadQueue.scala 152:68:@13028.4]
  wire  _T_15132; // @[LoadQueue.scala 151:92:@13030.4]
  wire  _T_15133; // @[LoadQueue.scala 152:41:@13031.4]
  wire  _T_15134; // @[LoadQueue.scala 153:30:@13032.4]
  wire  conflict_9_3; // @[LoadQueue.scala 152:68:@13033.4]
  wire  _T_15136; // @[LoadQueue.scala 151:92:@13035.4]
  wire  _T_15137; // @[LoadQueue.scala 152:41:@13036.4]
  wire  _T_15138; // @[LoadQueue.scala 153:30:@13037.4]
  wire  conflict_9_4; // @[LoadQueue.scala 152:68:@13038.4]
  wire  _T_15140; // @[LoadQueue.scala 151:92:@13040.4]
  wire  _T_15141; // @[LoadQueue.scala 152:41:@13041.4]
  wire  _T_15142; // @[LoadQueue.scala 153:30:@13042.4]
  wire  conflict_9_5; // @[LoadQueue.scala 152:68:@13043.4]
  wire  _T_15144; // @[LoadQueue.scala 151:92:@13045.4]
  wire  _T_15145; // @[LoadQueue.scala 152:41:@13046.4]
  wire  _T_15146; // @[LoadQueue.scala 153:30:@13047.4]
  wire  conflict_9_6; // @[LoadQueue.scala 152:68:@13048.4]
  wire  _T_15148; // @[LoadQueue.scala 151:92:@13050.4]
  wire  _T_15149; // @[LoadQueue.scala 152:41:@13051.4]
  wire  _T_15150; // @[LoadQueue.scala 153:30:@13052.4]
  wire  conflict_9_7; // @[LoadQueue.scala 152:68:@13053.4]
  wire  _T_15152; // @[LoadQueue.scala 151:92:@13055.4]
  wire  _T_15153; // @[LoadQueue.scala 152:41:@13056.4]
  wire  _T_15154; // @[LoadQueue.scala 153:30:@13057.4]
  wire  conflict_9_8; // @[LoadQueue.scala 152:68:@13058.4]
  wire  _T_15156; // @[LoadQueue.scala 151:92:@13060.4]
  wire  _T_15157; // @[LoadQueue.scala 152:41:@13061.4]
  wire  _T_15158; // @[LoadQueue.scala 153:30:@13062.4]
  wire  conflict_9_9; // @[LoadQueue.scala 152:68:@13063.4]
  wire  _T_15160; // @[LoadQueue.scala 151:92:@13065.4]
  wire  _T_15161; // @[LoadQueue.scala 152:41:@13066.4]
  wire  _T_15162; // @[LoadQueue.scala 153:30:@13067.4]
  wire  conflict_9_10; // @[LoadQueue.scala 152:68:@13068.4]
  wire  _T_15164; // @[LoadQueue.scala 151:92:@13070.4]
  wire  _T_15165; // @[LoadQueue.scala 152:41:@13071.4]
  wire  _T_15166; // @[LoadQueue.scala 153:30:@13072.4]
  wire  conflict_9_11; // @[LoadQueue.scala 152:68:@13073.4]
  wire  _T_15168; // @[LoadQueue.scala 151:92:@13075.4]
  wire  _T_15169; // @[LoadQueue.scala 152:41:@13076.4]
  wire  _T_15170; // @[LoadQueue.scala 153:30:@13077.4]
  wire  conflict_9_12; // @[LoadQueue.scala 152:68:@13078.4]
  wire  _T_15172; // @[LoadQueue.scala 151:92:@13080.4]
  wire  _T_15173; // @[LoadQueue.scala 152:41:@13081.4]
  wire  _T_15174; // @[LoadQueue.scala 153:30:@13082.4]
  wire  conflict_9_13; // @[LoadQueue.scala 152:68:@13083.4]
  wire  _T_15176; // @[LoadQueue.scala 151:92:@13085.4]
  wire  _T_15177; // @[LoadQueue.scala 152:41:@13086.4]
  wire  _T_15178; // @[LoadQueue.scala 153:30:@13087.4]
  wire  conflict_9_14; // @[LoadQueue.scala 152:68:@13088.4]
  wire  _T_15180; // @[LoadQueue.scala 151:92:@13090.4]
  wire  _T_15181; // @[LoadQueue.scala 152:41:@13091.4]
  wire  _T_15182; // @[LoadQueue.scala 153:30:@13092.4]
  wire  conflict_9_15; // @[LoadQueue.scala 152:68:@13093.4]
  wire  _T_15184; // @[LoadQueue.scala 151:92:@13095.4]
  wire  _T_15185; // @[LoadQueue.scala 152:41:@13096.4]
  wire  _T_15186; // @[LoadQueue.scala 153:30:@13097.4]
  wire  conflict_10_0; // @[LoadQueue.scala 152:68:@13098.4]
  wire  _T_15188; // @[LoadQueue.scala 151:92:@13100.4]
  wire  _T_15189; // @[LoadQueue.scala 152:41:@13101.4]
  wire  _T_15190; // @[LoadQueue.scala 153:30:@13102.4]
  wire  conflict_10_1; // @[LoadQueue.scala 152:68:@13103.4]
  wire  _T_15192; // @[LoadQueue.scala 151:92:@13105.4]
  wire  _T_15193; // @[LoadQueue.scala 152:41:@13106.4]
  wire  _T_15194; // @[LoadQueue.scala 153:30:@13107.4]
  wire  conflict_10_2; // @[LoadQueue.scala 152:68:@13108.4]
  wire  _T_15196; // @[LoadQueue.scala 151:92:@13110.4]
  wire  _T_15197; // @[LoadQueue.scala 152:41:@13111.4]
  wire  _T_15198; // @[LoadQueue.scala 153:30:@13112.4]
  wire  conflict_10_3; // @[LoadQueue.scala 152:68:@13113.4]
  wire  _T_15200; // @[LoadQueue.scala 151:92:@13115.4]
  wire  _T_15201; // @[LoadQueue.scala 152:41:@13116.4]
  wire  _T_15202; // @[LoadQueue.scala 153:30:@13117.4]
  wire  conflict_10_4; // @[LoadQueue.scala 152:68:@13118.4]
  wire  _T_15204; // @[LoadQueue.scala 151:92:@13120.4]
  wire  _T_15205; // @[LoadQueue.scala 152:41:@13121.4]
  wire  _T_15206; // @[LoadQueue.scala 153:30:@13122.4]
  wire  conflict_10_5; // @[LoadQueue.scala 152:68:@13123.4]
  wire  _T_15208; // @[LoadQueue.scala 151:92:@13125.4]
  wire  _T_15209; // @[LoadQueue.scala 152:41:@13126.4]
  wire  _T_15210; // @[LoadQueue.scala 153:30:@13127.4]
  wire  conflict_10_6; // @[LoadQueue.scala 152:68:@13128.4]
  wire  _T_15212; // @[LoadQueue.scala 151:92:@13130.4]
  wire  _T_15213; // @[LoadQueue.scala 152:41:@13131.4]
  wire  _T_15214; // @[LoadQueue.scala 153:30:@13132.4]
  wire  conflict_10_7; // @[LoadQueue.scala 152:68:@13133.4]
  wire  _T_15216; // @[LoadQueue.scala 151:92:@13135.4]
  wire  _T_15217; // @[LoadQueue.scala 152:41:@13136.4]
  wire  _T_15218; // @[LoadQueue.scala 153:30:@13137.4]
  wire  conflict_10_8; // @[LoadQueue.scala 152:68:@13138.4]
  wire  _T_15220; // @[LoadQueue.scala 151:92:@13140.4]
  wire  _T_15221; // @[LoadQueue.scala 152:41:@13141.4]
  wire  _T_15222; // @[LoadQueue.scala 153:30:@13142.4]
  wire  conflict_10_9; // @[LoadQueue.scala 152:68:@13143.4]
  wire  _T_15224; // @[LoadQueue.scala 151:92:@13145.4]
  wire  _T_15225; // @[LoadQueue.scala 152:41:@13146.4]
  wire  _T_15226; // @[LoadQueue.scala 153:30:@13147.4]
  wire  conflict_10_10; // @[LoadQueue.scala 152:68:@13148.4]
  wire  _T_15228; // @[LoadQueue.scala 151:92:@13150.4]
  wire  _T_15229; // @[LoadQueue.scala 152:41:@13151.4]
  wire  _T_15230; // @[LoadQueue.scala 153:30:@13152.4]
  wire  conflict_10_11; // @[LoadQueue.scala 152:68:@13153.4]
  wire  _T_15232; // @[LoadQueue.scala 151:92:@13155.4]
  wire  _T_15233; // @[LoadQueue.scala 152:41:@13156.4]
  wire  _T_15234; // @[LoadQueue.scala 153:30:@13157.4]
  wire  conflict_10_12; // @[LoadQueue.scala 152:68:@13158.4]
  wire  _T_15236; // @[LoadQueue.scala 151:92:@13160.4]
  wire  _T_15237; // @[LoadQueue.scala 152:41:@13161.4]
  wire  _T_15238; // @[LoadQueue.scala 153:30:@13162.4]
  wire  conflict_10_13; // @[LoadQueue.scala 152:68:@13163.4]
  wire  _T_15240; // @[LoadQueue.scala 151:92:@13165.4]
  wire  _T_15241; // @[LoadQueue.scala 152:41:@13166.4]
  wire  _T_15242; // @[LoadQueue.scala 153:30:@13167.4]
  wire  conflict_10_14; // @[LoadQueue.scala 152:68:@13168.4]
  wire  _T_15244; // @[LoadQueue.scala 151:92:@13170.4]
  wire  _T_15245; // @[LoadQueue.scala 152:41:@13171.4]
  wire  _T_15246; // @[LoadQueue.scala 153:30:@13172.4]
  wire  conflict_10_15; // @[LoadQueue.scala 152:68:@13173.4]
  wire  _T_15248; // @[LoadQueue.scala 151:92:@13175.4]
  wire  _T_15249; // @[LoadQueue.scala 152:41:@13176.4]
  wire  _T_15250; // @[LoadQueue.scala 153:30:@13177.4]
  wire  conflict_11_0; // @[LoadQueue.scala 152:68:@13178.4]
  wire  _T_15252; // @[LoadQueue.scala 151:92:@13180.4]
  wire  _T_15253; // @[LoadQueue.scala 152:41:@13181.4]
  wire  _T_15254; // @[LoadQueue.scala 153:30:@13182.4]
  wire  conflict_11_1; // @[LoadQueue.scala 152:68:@13183.4]
  wire  _T_15256; // @[LoadQueue.scala 151:92:@13185.4]
  wire  _T_15257; // @[LoadQueue.scala 152:41:@13186.4]
  wire  _T_15258; // @[LoadQueue.scala 153:30:@13187.4]
  wire  conflict_11_2; // @[LoadQueue.scala 152:68:@13188.4]
  wire  _T_15260; // @[LoadQueue.scala 151:92:@13190.4]
  wire  _T_15261; // @[LoadQueue.scala 152:41:@13191.4]
  wire  _T_15262; // @[LoadQueue.scala 153:30:@13192.4]
  wire  conflict_11_3; // @[LoadQueue.scala 152:68:@13193.4]
  wire  _T_15264; // @[LoadQueue.scala 151:92:@13195.4]
  wire  _T_15265; // @[LoadQueue.scala 152:41:@13196.4]
  wire  _T_15266; // @[LoadQueue.scala 153:30:@13197.4]
  wire  conflict_11_4; // @[LoadQueue.scala 152:68:@13198.4]
  wire  _T_15268; // @[LoadQueue.scala 151:92:@13200.4]
  wire  _T_15269; // @[LoadQueue.scala 152:41:@13201.4]
  wire  _T_15270; // @[LoadQueue.scala 153:30:@13202.4]
  wire  conflict_11_5; // @[LoadQueue.scala 152:68:@13203.4]
  wire  _T_15272; // @[LoadQueue.scala 151:92:@13205.4]
  wire  _T_15273; // @[LoadQueue.scala 152:41:@13206.4]
  wire  _T_15274; // @[LoadQueue.scala 153:30:@13207.4]
  wire  conflict_11_6; // @[LoadQueue.scala 152:68:@13208.4]
  wire  _T_15276; // @[LoadQueue.scala 151:92:@13210.4]
  wire  _T_15277; // @[LoadQueue.scala 152:41:@13211.4]
  wire  _T_15278; // @[LoadQueue.scala 153:30:@13212.4]
  wire  conflict_11_7; // @[LoadQueue.scala 152:68:@13213.4]
  wire  _T_15280; // @[LoadQueue.scala 151:92:@13215.4]
  wire  _T_15281; // @[LoadQueue.scala 152:41:@13216.4]
  wire  _T_15282; // @[LoadQueue.scala 153:30:@13217.4]
  wire  conflict_11_8; // @[LoadQueue.scala 152:68:@13218.4]
  wire  _T_15284; // @[LoadQueue.scala 151:92:@13220.4]
  wire  _T_15285; // @[LoadQueue.scala 152:41:@13221.4]
  wire  _T_15286; // @[LoadQueue.scala 153:30:@13222.4]
  wire  conflict_11_9; // @[LoadQueue.scala 152:68:@13223.4]
  wire  _T_15288; // @[LoadQueue.scala 151:92:@13225.4]
  wire  _T_15289; // @[LoadQueue.scala 152:41:@13226.4]
  wire  _T_15290; // @[LoadQueue.scala 153:30:@13227.4]
  wire  conflict_11_10; // @[LoadQueue.scala 152:68:@13228.4]
  wire  _T_15292; // @[LoadQueue.scala 151:92:@13230.4]
  wire  _T_15293; // @[LoadQueue.scala 152:41:@13231.4]
  wire  _T_15294; // @[LoadQueue.scala 153:30:@13232.4]
  wire  conflict_11_11; // @[LoadQueue.scala 152:68:@13233.4]
  wire  _T_15296; // @[LoadQueue.scala 151:92:@13235.4]
  wire  _T_15297; // @[LoadQueue.scala 152:41:@13236.4]
  wire  _T_15298; // @[LoadQueue.scala 153:30:@13237.4]
  wire  conflict_11_12; // @[LoadQueue.scala 152:68:@13238.4]
  wire  _T_15300; // @[LoadQueue.scala 151:92:@13240.4]
  wire  _T_15301; // @[LoadQueue.scala 152:41:@13241.4]
  wire  _T_15302; // @[LoadQueue.scala 153:30:@13242.4]
  wire  conflict_11_13; // @[LoadQueue.scala 152:68:@13243.4]
  wire  _T_15304; // @[LoadQueue.scala 151:92:@13245.4]
  wire  _T_15305; // @[LoadQueue.scala 152:41:@13246.4]
  wire  _T_15306; // @[LoadQueue.scala 153:30:@13247.4]
  wire  conflict_11_14; // @[LoadQueue.scala 152:68:@13248.4]
  wire  _T_15308; // @[LoadQueue.scala 151:92:@13250.4]
  wire  _T_15309; // @[LoadQueue.scala 152:41:@13251.4]
  wire  _T_15310; // @[LoadQueue.scala 153:30:@13252.4]
  wire  conflict_11_15; // @[LoadQueue.scala 152:68:@13253.4]
  wire  _T_15312; // @[LoadQueue.scala 151:92:@13255.4]
  wire  _T_15313; // @[LoadQueue.scala 152:41:@13256.4]
  wire  _T_15314; // @[LoadQueue.scala 153:30:@13257.4]
  wire  conflict_12_0; // @[LoadQueue.scala 152:68:@13258.4]
  wire  _T_15316; // @[LoadQueue.scala 151:92:@13260.4]
  wire  _T_15317; // @[LoadQueue.scala 152:41:@13261.4]
  wire  _T_15318; // @[LoadQueue.scala 153:30:@13262.4]
  wire  conflict_12_1; // @[LoadQueue.scala 152:68:@13263.4]
  wire  _T_15320; // @[LoadQueue.scala 151:92:@13265.4]
  wire  _T_15321; // @[LoadQueue.scala 152:41:@13266.4]
  wire  _T_15322; // @[LoadQueue.scala 153:30:@13267.4]
  wire  conflict_12_2; // @[LoadQueue.scala 152:68:@13268.4]
  wire  _T_15324; // @[LoadQueue.scala 151:92:@13270.4]
  wire  _T_15325; // @[LoadQueue.scala 152:41:@13271.4]
  wire  _T_15326; // @[LoadQueue.scala 153:30:@13272.4]
  wire  conflict_12_3; // @[LoadQueue.scala 152:68:@13273.4]
  wire  _T_15328; // @[LoadQueue.scala 151:92:@13275.4]
  wire  _T_15329; // @[LoadQueue.scala 152:41:@13276.4]
  wire  _T_15330; // @[LoadQueue.scala 153:30:@13277.4]
  wire  conflict_12_4; // @[LoadQueue.scala 152:68:@13278.4]
  wire  _T_15332; // @[LoadQueue.scala 151:92:@13280.4]
  wire  _T_15333; // @[LoadQueue.scala 152:41:@13281.4]
  wire  _T_15334; // @[LoadQueue.scala 153:30:@13282.4]
  wire  conflict_12_5; // @[LoadQueue.scala 152:68:@13283.4]
  wire  _T_15336; // @[LoadQueue.scala 151:92:@13285.4]
  wire  _T_15337; // @[LoadQueue.scala 152:41:@13286.4]
  wire  _T_15338; // @[LoadQueue.scala 153:30:@13287.4]
  wire  conflict_12_6; // @[LoadQueue.scala 152:68:@13288.4]
  wire  _T_15340; // @[LoadQueue.scala 151:92:@13290.4]
  wire  _T_15341; // @[LoadQueue.scala 152:41:@13291.4]
  wire  _T_15342; // @[LoadQueue.scala 153:30:@13292.4]
  wire  conflict_12_7; // @[LoadQueue.scala 152:68:@13293.4]
  wire  _T_15344; // @[LoadQueue.scala 151:92:@13295.4]
  wire  _T_15345; // @[LoadQueue.scala 152:41:@13296.4]
  wire  _T_15346; // @[LoadQueue.scala 153:30:@13297.4]
  wire  conflict_12_8; // @[LoadQueue.scala 152:68:@13298.4]
  wire  _T_15348; // @[LoadQueue.scala 151:92:@13300.4]
  wire  _T_15349; // @[LoadQueue.scala 152:41:@13301.4]
  wire  _T_15350; // @[LoadQueue.scala 153:30:@13302.4]
  wire  conflict_12_9; // @[LoadQueue.scala 152:68:@13303.4]
  wire  _T_15352; // @[LoadQueue.scala 151:92:@13305.4]
  wire  _T_15353; // @[LoadQueue.scala 152:41:@13306.4]
  wire  _T_15354; // @[LoadQueue.scala 153:30:@13307.4]
  wire  conflict_12_10; // @[LoadQueue.scala 152:68:@13308.4]
  wire  _T_15356; // @[LoadQueue.scala 151:92:@13310.4]
  wire  _T_15357; // @[LoadQueue.scala 152:41:@13311.4]
  wire  _T_15358; // @[LoadQueue.scala 153:30:@13312.4]
  wire  conflict_12_11; // @[LoadQueue.scala 152:68:@13313.4]
  wire  _T_15360; // @[LoadQueue.scala 151:92:@13315.4]
  wire  _T_15361; // @[LoadQueue.scala 152:41:@13316.4]
  wire  _T_15362; // @[LoadQueue.scala 153:30:@13317.4]
  wire  conflict_12_12; // @[LoadQueue.scala 152:68:@13318.4]
  wire  _T_15364; // @[LoadQueue.scala 151:92:@13320.4]
  wire  _T_15365; // @[LoadQueue.scala 152:41:@13321.4]
  wire  _T_15366; // @[LoadQueue.scala 153:30:@13322.4]
  wire  conflict_12_13; // @[LoadQueue.scala 152:68:@13323.4]
  wire  _T_15368; // @[LoadQueue.scala 151:92:@13325.4]
  wire  _T_15369; // @[LoadQueue.scala 152:41:@13326.4]
  wire  _T_15370; // @[LoadQueue.scala 153:30:@13327.4]
  wire  conflict_12_14; // @[LoadQueue.scala 152:68:@13328.4]
  wire  _T_15372; // @[LoadQueue.scala 151:92:@13330.4]
  wire  _T_15373; // @[LoadQueue.scala 152:41:@13331.4]
  wire  _T_15374; // @[LoadQueue.scala 153:30:@13332.4]
  wire  conflict_12_15; // @[LoadQueue.scala 152:68:@13333.4]
  wire  _T_15376; // @[LoadQueue.scala 151:92:@13335.4]
  wire  _T_15377; // @[LoadQueue.scala 152:41:@13336.4]
  wire  _T_15378; // @[LoadQueue.scala 153:30:@13337.4]
  wire  conflict_13_0; // @[LoadQueue.scala 152:68:@13338.4]
  wire  _T_15380; // @[LoadQueue.scala 151:92:@13340.4]
  wire  _T_15381; // @[LoadQueue.scala 152:41:@13341.4]
  wire  _T_15382; // @[LoadQueue.scala 153:30:@13342.4]
  wire  conflict_13_1; // @[LoadQueue.scala 152:68:@13343.4]
  wire  _T_15384; // @[LoadQueue.scala 151:92:@13345.4]
  wire  _T_15385; // @[LoadQueue.scala 152:41:@13346.4]
  wire  _T_15386; // @[LoadQueue.scala 153:30:@13347.4]
  wire  conflict_13_2; // @[LoadQueue.scala 152:68:@13348.4]
  wire  _T_15388; // @[LoadQueue.scala 151:92:@13350.4]
  wire  _T_15389; // @[LoadQueue.scala 152:41:@13351.4]
  wire  _T_15390; // @[LoadQueue.scala 153:30:@13352.4]
  wire  conflict_13_3; // @[LoadQueue.scala 152:68:@13353.4]
  wire  _T_15392; // @[LoadQueue.scala 151:92:@13355.4]
  wire  _T_15393; // @[LoadQueue.scala 152:41:@13356.4]
  wire  _T_15394; // @[LoadQueue.scala 153:30:@13357.4]
  wire  conflict_13_4; // @[LoadQueue.scala 152:68:@13358.4]
  wire  _T_15396; // @[LoadQueue.scala 151:92:@13360.4]
  wire  _T_15397; // @[LoadQueue.scala 152:41:@13361.4]
  wire  _T_15398; // @[LoadQueue.scala 153:30:@13362.4]
  wire  conflict_13_5; // @[LoadQueue.scala 152:68:@13363.4]
  wire  _T_15400; // @[LoadQueue.scala 151:92:@13365.4]
  wire  _T_15401; // @[LoadQueue.scala 152:41:@13366.4]
  wire  _T_15402; // @[LoadQueue.scala 153:30:@13367.4]
  wire  conflict_13_6; // @[LoadQueue.scala 152:68:@13368.4]
  wire  _T_15404; // @[LoadQueue.scala 151:92:@13370.4]
  wire  _T_15405; // @[LoadQueue.scala 152:41:@13371.4]
  wire  _T_15406; // @[LoadQueue.scala 153:30:@13372.4]
  wire  conflict_13_7; // @[LoadQueue.scala 152:68:@13373.4]
  wire  _T_15408; // @[LoadQueue.scala 151:92:@13375.4]
  wire  _T_15409; // @[LoadQueue.scala 152:41:@13376.4]
  wire  _T_15410; // @[LoadQueue.scala 153:30:@13377.4]
  wire  conflict_13_8; // @[LoadQueue.scala 152:68:@13378.4]
  wire  _T_15412; // @[LoadQueue.scala 151:92:@13380.4]
  wire  _T_15413; // @[LoadQueue.scala 152:41:@13381.4]
  wire  _T_15414; // @[LoadQueue.scala 153:30:@13382.4]
  wire  conflict_13_9; // @[LoadQueue.scala 152:68:@13383.4]
  wire  _T_15416; // @[LoadQueue.scala 151:92:@13385.4]
  wire  _T_15417; // @[LoadQueue.scala 152:41:@13386.4]
  wire  _T_15418; // @[LoadQueue.scala 153:30:@13387.4]
  wire  conflict_13_10; // @[LoadQueue.scala 152:68:@13388.4]
  wire  _T_15420; // @[LoadQueue.scala 151:92:@13390.4]
  wire  _T_15421; // @[LoadQueue.scala 152:41:@13391.4]
  wire  _T_15422; // @[LoadQueue.scala 153:30:@13392.4]
  wire  conflict_13_11; // @[LoadQueue.scala 152:68:@13393.4]
  wire  _T_15424; // @[LoadQueue.scala 151:92:@13395.4]
  wire  _T_15425; // @[LoadQueue.scala 152:41:@13396.4]
  wire  _T_15426; // @[LoadQueue.scala 153:30:@13397.4]
  wire  conflict_13_12; // @[LoadQueue.scala 152:68:@13398.4]
  wire  _T_15428; // @[LoadQueue.scala 151:92:@13400.4]
  wire  _T_15429; // @[LoadQueue.scala 152:41:@13401.4]
  wire  _T_15430; // @[LoadQueue.scala 153:30:@13402.4]
  wire  conflict_13_13; // @[LoadQueue.scala 152:68:@13403.4]
  wire  _T_15432; // @[LoadQueue.scala 151:92:@13405.4]
  wire  _T_15433; // @[LoadQueue.scala 152:41:@13406.4]
  wire  _T_15434; // @[LoadQueue.scala 153:30:@13407.4]
  wire  conflict_13_14; // @[LoadQueue.scala 152:68:@13408.4]
  wire  _T_15436; // @[LoadQueue.scala 151:92:@13410.4]
  wire  _T_15437; // @[LoadQueue.scala 152:41:@13411.4]
  wire  _T_15438; // @[LoadQueue.scala 153:30:@13412.4]
  wire  conflict_13_15; // @[LoadQueue.scala 152:68:@13413.4]
  wire  _T_15440; // @[LoadQueue.scala 151:92:@13415.4]
  wire  _T_15441; // @[LoadQueue.scala 152:41:@13416.4]
  wire  _T_15442; // @[LoadQueue.scala 153:30:@13417.4]
  wire  conflict_14_0; // @[LoadQueue.scala 152:68:@13418.4]
  wire  _T_15444; // @[LoadQueue.scala 151:92:@13420.4]
  wire  _T_15445; // @[LoadQueue.scala 152:41:@13421.4]
  wire  _T_15446; // @[LoadQueue.scala 153:30:@13422.4]
  wire  conflict_14_1; // @[LoadQueue.scala 152:68:@13423.4]
  wire  _T_15448; // @[LoadQueue.scala 151:92:@13425.4]
  wire  _T_15449; // @[LoadQueue.scala 152:41:@13426.4]
  wire  _T_15450; // @[LoadQueue.scala 153:30:@13427.4]
  wire  conflict_14_2; // @[LoadQueue.scala 152:68:@13428.4]
  wire  _T_15452; // @[LoadQueue.scala 151:92:@13430.4]
  wire  _T_15453; // @[LoadQueue.scala 152:41:@13431.4]
  wire  _T_15454; // @[LoadQueue.scala 153:30:@13432.4]
  wire  conflict_14_3; // @[LoadQueue.scala 152:68:@13433.4]
  wire  _T_15456; // @[LoadQueue.scala 151:92:@13435.4]
  wire  _T_15457; // @[LoadQueue.scala 152:41:@13436.4]
  wire  _T_15458; // @[LoadQueue.scala 153:30:@13437.4]
  wire  conflict_14_4; // @[LoadQueue.scala 152:68:@13438.4]
  wire  _T_15460; // @[LoadQueue.scala 151:92:@13440.4]
  wire  _T_15461; // @[LoadQueue.scala 152:41:@13441.4]
  wire  _T_15462; // @[LoadQueue.scala 153:30:@13442.4]
  wire  conflict_14_5; // @[LoadQueue.scala 152:68:@13443.4]
  wire  _T_15464; // @[LoadQueue.scala 151:92:@13445.4]
  wire  _T_15465; // @[LoadQueue.scala 152:41:@13446.4]
  wire  _T_15466; // @[LoadQueue.scala 153:30:@13447.4]
  wire  conflict_14_6; // @[LoadQueue.scala 152:68:@13448.4]
  wire  _T_15468; // @[LoadQueue.scala 151:92:@13450.4]
  wire  _T_15469; // @[LoadQueue.scala 152:41:@13451.4]
  wire  _T_15470; // @[LoadQueue.scala 153:30:@13452.4]
  wire  conflict_14_7; // @[LoadQueue.scala 152:68:@13453.4]
  wire  _T_15472; // @[LoadQueue.scala 151:92:@13455.4]
  wire  _T_15473; // @[LoadQueue.scala 152:41:@13456.4]
  wire  _T_15474; // @[LoadQueue.scala 153:30:@13457.4]
  wire  conflict_14_8; // @[LoadQueue.scala 152:68:@13458.4]
  wire  _T_15476; // @[LoadQueue.scala 151:92:@13460.4]
  wire  _T_15477; // @[LoadQueue.scala 152:41:@13461.4]
  wire  _T_15478; // @[LoadQueue.scala 153:30:@13462.4]
  wire  conflict_14_9; // @[LoadQueue.scala 152:68:@13463.4]
  wire  _T_15480; // @[LoadQueue.scala 151:92:@13465.4]
  wire  _T_15481; // @[LoadQueue.scala 152:41:@13466.4]
  wire  _T_15482; // @[LoadQueue.scala 153:30:@13467.4]
  wire  conflict_14_10; // @[LoadQueue.scala 152:68:@13468.4]
  wire  _T_15484; // @[LoadQueue.scala 151:92:@13470.4]
  wire  _T_15485; // @[LoadQueue.scala 152:41:@13471.4]
  wire  _T_15486; // @[LoadQueue.scala 153:30:@13472.4]
  wire  conflict_14_11; // @[LoadQueue.scala 152:68:@13473.4]
  wire  _T_15488; // @[LoadQueue.scala 151:92:@13475.4]
  wire  _T_15489; // @[LoadQueue.scala 152:41:@13476.4]
  wire  _T_15490; // @[LoadQueue.scala 153:30:@13477.4]
  wire  conflict_14_12; // @[LoadQueue.scala 152:68:@13478.4]
  wire  _T_15492; // @[LoadQueue.scala 151:92:@13480.4]
  wire  _T_15493; // @[LoadQueue.scala 152:41:@13481.4]
  wire  _T_15494; // @[LoadQueue.scala 153:30:@13482.4]
  wire  conflict_14_13; // @[LoadQueue.scala 152:68:@13483.4]
  wire  _T_15496; // @[LoadQueue.scala 151:92:@13485.4]
  wire  _T_15497; // @[LoadQueue.scala 152:41:@13486.4]
  wire  _T_15498; // @[LoadQueue.scala 153:30:@13487.4]
  wire  conflict_14_14; // @[LoadQueue.scala 152:68:@13488.4]
  wire  _T_15500; // @[LoadQueue.scala 151:92:@13490.4]
  wire  _T_15501; // @[LoadQueue.scala 152:41:@13491.4]
  wire  _T_15502; // @[LoadQueue.scala 153:30:@13492.4]
  wire  conflict_14_15; // @[LoadQueue.scala 152:68:@13493.4]
  wire  _T_15504; // @[LoadQueue.scala 151:92:@13495.4]
  wire  _T_15505; // @[LoadQueue.scala 152:41:@13496.4]
  wire  _T_15506; // @[LoadQueue.scala 153:30:@13497.4]
  wire  conflict_15_0; // @[LoadQueue.scala 152:68:@13498.4]
  wire  _T_15508; // @[LoadQueue.scala 151:92:@13500.4]
  wire  _T_15509; // @[LoadQueue.scala 152:41:@13501.4]
  wire  _T_15510; // @[LoadQueue.scala 153:30:@13502.4]
  wire  conflict_15_1; // @[LoadQueue.scala 152:68:@13503.4]
  wire  _T_15512; // @[LoadQueue.scala 151:92:@13505.4]
  wire  _T_15513; // @[LoadQueue.scala 152:41:@13506.4]
  wire  _T_15514; // @[LoadQueue.scala 153:30:@13507.4]
  wire  conflict_15_2; // @[LoadQueue.scala 152:68:@13508.4]
  wire  _T_15516; // @[LoadQueue.scala 151:92:@13510.4]
  wire  _T_15517; // @[LoadQueue.scala 152:41:@13511.4]
  wire  _T_15518; // @[LoadQueue.scala 153:30:@13512.4]
  wire  conflict_15_3; // @[LoadQueue.scala 152:68:@13513.4]
  wire  _T_15520; // @[LoadQueue.scala 151:92:@13515.4]
  wire  _T_15521; // @[LoadQueue.scala 152:41:@13516.4]
  wire  _T_15522; // @[LoadQueue.scala 153:30:@13517.4]
  wire  conflict_15_4; // @[LoadQueue.scala 152:68:@13518.4]
  wire  _T_15524; // @[LoadQueue.scala 151:92:@13520.4]
  wire  _T_15525; // @[LoadQueue.scala 152:41:@13521.4]
  wire  _T_15526; // @[LoadQueue.scala 153:30:@13522.4]
  wire  conflict_15_5; // @[LoadQueue.scala 152:68:@13523.4]
  wire  _T_15528; // @[LoadQueue.scala 151:92:@13525.4]
  wire  _T_15529; // @[LoadQueue.scala 152:41:@13526.4]
  wire  _T_15530; // @[LoadQueue.scala 153:30:@13527.4]
  wire  conflict_15_6; // @[LoadQueue.scala 152:68:@13528.4]
  wire  _T_15532; // @[LoadQueue.scala 151:92:@13530.4]
  wire  _T_15533; // @[LoadQueue.scala 152:41:@13531.4]
  wire  _T_15534; // @[LoadQueue.scala 153:30:@13532.4]
  wire  conflict_15_7; // @[LoadQueue.scala 152:68:@13533.4]
  wire  _T_15536; // @[LoadQueue.scala 151:92:@13535.4]
  wire  _T_15537; // @[LoadQueue.scala 152:41:@13536.4]
  wire  _T_15538; // @[LoadQueue.scala 153:30:@13537.4]
  wire  conflict_15_8; // @[LoadQueue.scala 152:68:@13538.4]
  wire  _T_15540; // @[LoadQueue.scala 151:92:@13540.4]
  wire  _T_15541; // @[LoadQueue.scala 152:41:@13541.4]
  wire  _T_15542; // @[LoadQueue.scala 153:30:@13542.4]
  wire  conflict_15_9; // @[LoadQueue.scala 152:68:@13543.4]
  wire  _T_15544; // @[LoadQueue.scala 151:92:@13545.4]
  wire  _T_15545; // @[LoadQueue.scala 152:41:@13546.4]
  wire  _T_15546; // @[LoadQueue.scala 153:30:@13547.4]
  wire  conflict_15_10; // @[LoadQueue.scala 152:68:@13548.4]
  wire  _T_15548; // @[LoadQueue.scala 151:92:@13550.4]
  wire  _T_15549; // @[LoadQueue.scala 152:41:@13551.4]
  wire  _T_15550; // @[LoadQueue.scala 153:30:@13552.4]
  wire  conflict_15_11; // @[LoadQueue.scala 152:68:@13553.4]
  wire  _T_15552; // @[LoadQueue.scala 151:92:@13555.4]
  wire  _T_15553; // @[LoadQueue.scala 152:41:@13556.4]
  wire  _T_15554; // @[LoadQueue.scala 153:30:@13557.4]
  wire  conflict_15_12; // @[LoadQueue.scala 152:68:@13558.4]
  wire  _T_15556; // @[LoadQueue.scala 151:92:@13560.4]
  wire  _T_15557; // @[LoadQueue.scala 152:41:@13561.4]
  wire  _T_15558; // @[LoadQueue.scala 153:30:@13562.4]
  wire  conflict_15_13; // @[LoadQueue.scala 152:68:@13563.4]
  wire  _T_15560; // @[LoadQueue.scala 151:92:@13565.4]
  wire  _T_15561; // @[LoadQueue.scala 152:41:@13566.4]
  wire  _T_15562; // @[LoadQueue.scala 153:30:@13567.4]
  wire  conflict_15_14; // @[LoadQueue.scala 152:68:@13568.4]
  wire  _T_15564; // @[LoadQueue.scala 151:92:@13570.4]
  wire  _T_15565; // @[LoadQueue.scala 152:41:@13571.4]
  wire  _T_15566; // @[LoadQueue.scala 153:30:@13572.4]
  wire  conflict_15_15; // @[LoadQueue.scala 152:68:@13573.4]
  wire  _T_16799; // @[LoadQueue.scala 163:13:@13576.4]
  wire  storeAddrNotKnownFlags_0_0; // @[LoadQueue.scala 163:19:@13577.4]
  wire  _T_16802; // @[LoadQueue.scala 163:13:@13578.4]
  wire  storeAddrNotKnownFlags_0_1; // @[LoadQueue.scala 163:19:@13579.4]
  wire  _T_16805; // @[LoadQueue.scala 163:13:@13580.4]
  wire  storeAddrNotKnownFlags_0_2; // @[LoadQueue.scala 163:19:@13581.4]
  wire  _T_16808; // @[LoadQueue.scala 163:13:@13582.4]
  wire  storeAddrNotKnownFlags_0_3; // @[LoadQueue.scala 163:19:@13583.4]
  wire  _T_16811; // @[LoadQueue.scala 163:13:@13584.4]
  wire  storeAddrNotKnownFlags_0_4; // @[LoadQueue.scala 163:19:@13585.4]
  wire  _T_16814; // @[LoadQueue.scala 163:13:@13586.4]
  wire  storeAddrNotKnownFlags_0_5; // @[LoadQueue.scala 163:19:@13587.4]
  wire  _T_16817; // @[LoadQueue.scala 163:13:@13588.4]
  wire  storeAddrNotKnownFlags_0_6; // @[LoadQueue.scala 163:19:@13589.4]
  wire  _T_16820; // @[LoadQueue.scala 163:13:@13590.4]
  wire  storeAddrNotKnownFlags_0_7; // @[LoadQueue.scala 163:19:@13591.4]
  wire  _T_16823; // @[LoadQueue.scala 163:13:@13592.4]
  wire  storeAddrNotKnownFlags_0_8; // @[LoadQueue.scala 163:19:@13593.4]
  wire  _T_16826; // @[LoadQueue.scala 163:13:@13594.4]
  wire  storeAddrNotKnownFlags_0_9; // @[LoadQueue.scala 163:19:@13595.4]
  wire  _T_16829; // @[LoadQueue.scala 163:13:@13596.4]
  wire  storeAddrNotKnownFlags_0_10; // @[LoadQueue.scala 163:19:@13597.4]
  wire  _T_16832; // @[LoadQueue.scala 163:13:@13598.4]
  wire  storeAddrNotKnownFlags_0_11; // @[LoadQueue.scala 163:19:@13599.4]
  wire  _T_16835; // @[LoadQueue.scala 163:13:@13600.4]
  wire  storeAddrNotKnownFlags_0_12; // @[LoadQueue.scala 163:19:@13601.4]
  wire  _T_16838; // @[LoadQueue.scala 163:13:@13602.4]
  wire  storeAddrNotKnownFlags_0_13; // @[LoadQueue.scala 163:19:@13603.4]
  wire  _T_16841; // @[LoadQueue.scala 163:13:@13604.4]
  wire  storeAddrNotKnownFlags_0_14; // @[LoadQueue.scala 163:19:@13605.4]
  wire  _T_16844; // @[LoadQueue.scala 163:13:@13606.4]
  wire  storeAddrNotKnownFlags_0_15; // @[LoadQueue.scala 163:19:@13607.4]
  wire  storeAddrNotKnownFlags_1_0; // @[LoadQueue.scala 163:19:@13625.4]
  wire  storeAddrNotKnownFlags_1_1; // @[LoadQueue.scala 163:19:@13627.4]
  wire  storeAddrNotKnownFlags_1_2; // @[LoadQueue.scala 163:19:@13629.4]
  wire  storeAddrNotKnownFlags_1_3; // @[LoadQueue.scala 163:19:@13631.4]
  wire  storeAddrNotKnownFlags_1_4; // @[LoadQueue.scala 163:19:@13633.4]
  wire  storeAddrNotKnownFlags_1_5; // @[LoadQueue.scala 163:19:@13635.4]
  wire  storeAddrNotKnownFlags_1_6; // @[LoadQueue.scala 163:19:@13637.4]
  wire  storeAddrNotKnownFlags_1_7; // @[LoadQueue.scala 163:19:@13639.4]
  wire  storeAddrNotKnownFlags_1_8; // @[LoadQueue.scala 163:19:@13641.4]
  wire  storeAddrNotKnownFlags_1_9; // @[LoadQueue.scala 163:19:@13643.4]
  wire  storeAddrNotKnownFlags_1_10; // @[LoadQueue.scala 163:19:@13645.4]
  wire  storeAddrNotKnownFlags_1_11; // @[LoadQueue.scala 163:19:@13647.4]
  wire  storeAddrNotKnownFlags_1_12; // @[LoadQueue.scala 163:19:@13649.4]
  wire  storeAddrNotKnownFlags_1_13; // @[LoadQueue.scala 163:19:@13651.4]
  wire  storeAddrNotKnownFlags_1_14; // @[LoadQueue.scala 163:19:@13653.4]
  wire  storeAddrNotKnownFlags_1_15; // @[LoadQueue.scala 163:19:@13655.4]
  wire  storeAddrNotKnownFlags_2_0; // @[LoadQueue.scala 163:19:@13673.4]
  wire  storeAddrNotKnownFlags_2_1; // @[LoadQueue.scala 163:19:@13675.4]
  wire  storeAddrNotKnownFlags_2_2; // @[LoadQueue.scala 163:19:@13677.4]
  wire  storeAddrNotKnownFlags_2_3; // @[LoadQueue.scala 163:19:@13679.4]
  wire  storeAddrNotKnownFlags_2_4; // @[LoadQueue.scala 163:19:@13681.4]
  wire  storeAddrNotKnownFlags_2_5; // @[LoadQueue.scala 163:19:@13683.4]
  wire  storeAddrNotKnownFlags_2_6; // @[LoadQueue.scala 163:19:@13685.4]
  wire  storeAddrNotKnownFlags_2_7; // @[LoadQueue.scala 163:19:@13687.4]
  wire  storeAddrNotKnownFlags_2_8; // @[LoadQueue.scala 163:19:@13689.4]
  wire  storeAddrNotKnownFlags_2_9; // @[LoadQueue.scala 163:19:@13691.4]
  wire  storeAddrNotKnownFlags_2_10; // @[LoadQueue.scala 163:19:@13693.4]
  wire  storeAddrNotKnownFlags_2_11; // @[LoadQueue.scala 163:19:@13695.4]
  wire  storeAddrNotKnownFlags_2_12; // @[LoadQueue.scala 163:19:@13697.4]
  wire  storeAddrNotKnownFlags_2_13; // @[LoadQueue.scala 163:19:@13699.4]
  wire  storeAddrNotKnownFlags_2_14; // @[LoadQueue.scala 163:19:@13701.4]
  wire  storeAddrNotKnownFlags_2_15; // @[LoadQueue.scala 163:19:@13703.4]
  wire  storeAddrNotKnownFlags_3_0; // @[LoadQueue.scala 163:19:@13721.4]
  wire  storeAddrNotKnownFlags_3_1; // @[LoadQueue.scala 163:19:@13723.4]
  wire  storeAddrNotKnownFlags_3_2; // @[LoadQueue.scala 163:19:@13725.4]
  wire  storeAddrNotKnownFlags_3_3; // @[LoadQueue.scala 163:19:@13727.4]
  wire  storeAddrNotKnownFlags_3_4; // @[LoadQueue.scala 163:19:@13729.4]
  wire  storeAddrNotKnownFlags_3_5; // @[LoadQueue.scala 163:19:@13731.4]
  wire  storeAddrNotKnownFlags_3_6; // @[LoadQueue.scala 163:19:@13733.4]
  wire  storeAddrNotKnownFlags_3_7; // @[LoadQueue.scala 163:19:@13735.4]
  wire  storeAddrNotKnownFlags_3_8; // @[LoadQueue.scala 163:19:@13737.4]
  wire  storeAddrNotKnownFlags_3_9; // @[LoadQueue.scala 163:19:@13739.4]
  wire  storeAddrNotKnownFlags_3_10; // @[LoadQueue.scala 163:19:@13741.4]
  wire  storeAddrNotKnownFlags_3_11; // @[LoadQueue.scala 163:19:@13743.4]
  wire  storeAddrNotKnownFlags_3_12; // @[LoadQueue.scala 163:19:@13745.4]
  wire  storeAddrNotKnownFlags_3_13; // @[LoadQueue.scala 163:19:@13747.4]
  wire  storeAddrNotKnownFlags_3_14; // @[LoadQueue.scala 163:19:@13749.4]
  wire  storeAddrNotKnownFlags_3_15; // @[LoadQueue.scala 163:19:@13751.4]
  wire  storeAddrNotKnownFlags_4_0; // @[LoadQueue.scala 163:19:@13769.4]
  wire  storeAddrNotKnownFlags_4_1; // @[LoadQueue.scala 163:19:@13771.4]
  wire  storeAddrNotKnownFlags_4_2; // @[LoadQueue.scala 163:19:@13773.4]
  wire  storeAddrNotKnownFlags_4_3; // @[LoadQueue.scala 163:19:@13775.4]
  wire  storeAddrNotKnownFlags_4_4; // @[LoadQueue.scala 163:19:@13777.4]
  wire  storeAddrNotKnownFlags_4_5; // @[LoadQueue.scala 163:19:@13779.4]
  wire  storeAddrNotKnownFlags_4_6; // @[LoadQueue.scala 163:19:@13781.4]
  wire  storeAddrNotKnownFlags_4_7; // @[LoadQueue.scala 163:19:@13783.4]
  wire  storeAddrNotKnownFlags_4_8; // @[LoadQueue.scala 163:19:@13785.4]
  wire  storeAddrNotKnownFlags_4_9; // @[LoadQueue.scala 163:19:@13787.4]
  wire  storeAddrNotKnownFlags_4_10; // @[LoadQueue.scala 163:19:@13789.4]
  wire  storeAddrNotKnownFlags_4_11; // @[LoadQueue.scala 163:19:@13791.4]
  wire  storeAddrNotKnownFlags_4_12; // @[LoadQueue.scala 163:19:@13793.4]
  wire  storeAddrNotKnownFlags_4_13; // @[LoadQueue.scala 163:19:@13795.4]
  wire  storeAddrNotKnownFlags_4_14; // @[LoadQueue.scala 163:19:@13797.4]
  wire  storeAddrNotKnownFlags_4_15; // @[LoadQueue.scala 163:19:@13799.4]
  wire  storeAddrNotKnownFlags_5_0; // @[LoadQueue.scala 163:19:@13817.4]
  wire  storeAddrNotKnownFlags_5_1; // @[LoadQueue.scala 163:19:@13819.4]
  wire  storeAddrNotKnownFlags_5_2; // @[LoadQueue.scala 163:19:@13821.4]
  wire  storeAddrNotKnownFlags_5_3; // @[LoadQueue.scala 163:19:@13823.4]
  wire  storeAddrNotKnownFlags_5_4; // @[LoadQueue.scala 163:19:@13825.4]
  wire  storeAddrNotKnownFlags_5_5; // @[LoadQueue.scala 163:19:@13827.4]
  wire  storeAddrNotKnownFlags_5_6; // @[LoadQueue.scala 163:19:@13829.4]
  wire  storeAddrNotKnownFlags_5_7; // @[LoadQueue.scala 163:19:@13831.4]
  wire  storeAddrNotKnownFlags_5_8; // @[LoadQueue.scala 163:19:@13833.4]
  wire  storeAddrNotKnownFlags_5_9; // @[LoadQueue.scala 163:19:@13835.4]
  wire  storeAddrNotKnownFlags_5_10; // @[LoadQueue.scala 163:19:@13837.4]
  wire  storeAddrNotKnownFlags_5_11; // @[LoadQueue.scala 163:19:@13839.4]
  wire  storeAddrNotKnownFlags_5_12; // @[LoadQueue.scala 163:19:@13841.4]
  wire  storeAddrNotKnownFlags_5_13; // @[LoadQueue.scala 163:19:@13843.4]
  wire  storeAddrNotKnownFlags_5_14; // @[LoadQueue.scala 163:19:@13845.4]
  wire  storeAddrNotKnownFlags_5_15; // @[LoadQueue.scala 163:19:@13847.4]
  wire  storeAddrNotKnownFlags_6_0; // @[LoadQueue.scala 163:19:@13865.4]
  wire  storeAddrNotKnownFlags_6_1; // @[LoadQueue.scala 163:19:@13867.4]
  wire  storeAddrNotKnownFlags_6_2; // @[LoadQueue.scala 163:19:@13869.4]
  wire  storeAddrNotKnownFlags_6_3; // @[LoadQueue.scala 163:19:@13871.4]
  wire  storeAddrNotKnownFlags_6_4; // @[LoadQueue.scala 163:19:@13873.4]
  wire  storeAddrNotKnownFlags_6_5; // @[LoadQueue.scala 163:19:@13875.4]
  wire  storeAddrNotKnownFlags_6_6; // @[LoadQueue.scala 163:19:@13877.4]
  wire  storeAddrNotKnownFlags_6_7; // @[LoadQueue.scala 163:19:@13879.4]
  wire  storeAddrNotKnownFlags_6_8; // @[LoadQueue.scala 163:19:@13881.4]
  wire  storeAddrNotKnownFlags_6_9; // @[LoadQueue.scala 163:19:@13883.4]
  wire  storeAddrNotKnownFlags_6_10; // @[LoadQueue.scala 163:19:@13885.4]
  wire  storeAddrNotKnownFlags_6_11; // @[LoadQueue.scala 163:19:@13887.4]
  wire  storeAddrNotKnownFlags_6_12; // @[LoadQueue.scala 163:19:@13889.4]
  wire  storeAddrNotKnownFlags_6_13; // @[LoadQueue.scala 163:19:@13891.4]
  wire  storeAddrNotKnownFlags_6_14; // @[LoadQueue.scala 163:19:@13893.4]
  wire  storeAddrNotKnownFlags_6_15; // @[LoadQueue.scala 163:19:@13895.4]
  wire  storeAddrNotKnownFlags_7_0; // @[LoadQueue.scala 163:19:@13913.4]
  wire  storeAddrNotKnownFlags_7_1; // @[LoadQueue.scala 163:19:@13915.4]
  wire  storeAddrNotKnownFlags_7_2; // @[LoadQueue.scala 163:19:@13917.4]
  wire  storeAddrNotKnownFlags_7_3; // @[LoadQueue.scala 163:19:@13919.4]
  wire  storeAddrNotKnownFlags_7_4; // @[LoadQueue.scala 163:19:@13921.4]
  wire  storeAddrNotKnownFlags_7_5; // @[LoadQueue.scala 163:19:@13923.4]
  wire  storeAddrNotKnownFlags_7_6; // @[LoadQueue.scala 163:19:@13925.4]
  wire  storeAddrNotKnownFlags_7_7; // @[LoadQueue.scala 163:19:@13927.4]
  wire  storeAddrNotKnownFlags_7_8; // @[LoadQueue.scala 163:19:@13929.4]
  wire  storeAddrNotKnownFlags_7_9; // @[LoadQueue.scala 163:19:@13931.4]
  wire  storeAddrNotKnownFlags_7_10; // @[LoadQueue.scala 163:19:@13933.4]
  wire  storeAddrNotKnownFlags_7_11; // @[LoadQueue.scala 163:19:@13935.4]
  wire  storeAddrNotKnownFlags_7_12; // @[LoadQueue.scala 163:19:@13937.4]
  wire  storeAddrNotKnownFlags_7_13; // @[LoadQueue.scala 163:19:@13939.4]
  wire  storeAddrNotKnownFlags_7_14; // @[LoadQueue.scala 163:19:@13941.4]
  wire  storeAddrNotKnownFlags_7_15; // @[LoadQueue.scala 163:19:@13943.4]
  wire  storeAddrNotKnownFlags_8_0; // @[LoadQueue.scala 163:19:@13961.4]
  wire  storeAddrNotKnownFlags_8_1; // @[LoadQueue.scala 163:19:@13963.4]
  wire  storeAddrNotKnownFlags_8_2; // @[LoadQueue.scala 163:19:@13965.4]
  wire  storeAddrNotKnownFlags_8_3; // @[LoadQueue.scala 163:19:@13967.4]
  wire  storeAddrNotKnownFlags_8_4; // @[LoadQueue.scala 163:19:@13969.4]
  wire  storeAddrNotKnownFlags_8_5; // @[LoadQueue.scala 163:19:@13971.4]
  wire  storeAddrNotKnownFlags_8_6; // @[LoadQueue.scala 163:19:@13973.4]
  wire  storeAddrNotKnownFlags_8_7; // @[LoadQueue.scala 163:19:@13975.4]
  wire  storeAddrNotKnownFlags_8_8; // @[LoadQueue.scala 163:19:@13977.4]
  wire  storeAddrNotKnownFlags_8_9; // @[LoadQueue.scala 163:19:@13979.4]
  wire  storeAddrNotKnownFlags_8_10; // @[LoadQueue.scala 163:19:@13981.4]
  wire  storeAddrNotKnownFlags_8_11; // @[LoadQueue.scala 163:19:@13983.4]
  wire  storeAddrNotKnownFlags_8_12; // @[LoadQueue.scala 163:19:@13985.4]
  wire  storeAddrNotKnownFlags_8_13; // @[LoadQueue.scala 163:19:@13987.4]
  wire  storeAddrNotKnownFlags_8_14; // @[LoadQueue.scala 163:19:@13989.4]
  wire  storeAddrNotKnownFlags_8_15; // @[LoadQueue.scala 163:19:@13991.4]
  wire  storeAddrNotKnownFlags_9_0; // @[LoadQueue.scala 163:19:@14009.4]
  wire  storeAddrNotKnownFlags_9_1; // @[LoadQueue.scala 163:19:@14011.4]
  wire  storeAddrNotKnownFlags_9_2; // @[LoadQueue.scala 163:19:@14013.4]
  wire  storeAddrNotKnownFlags_9_3; // @[LoadQueue.scala 163:19:@14015.4]
  wire  storeAddrNotKnownFlags_9_4; // @[LoadQueue.scala 163:19:@14017.4]
  wire  storeAddrNotKnownFlags_9_5; // @[LoadQueue.scala 163:19:@14019.4]
  wire  storeAddrNotKnownFlags_9_6; // @[LoadQueue.scala 163:19:@14021.4]
  wire  storeAddrNotKnownFlags_9_7; // @[LoadQueue.scala 163:19:@14023.4]
  wire  storeAddrNotKnownFlags_9_8; // @[LoadQueue.scala 163:19:@14025.4]
  wire  storeAddrNotKnownFlags_9_9; // @[LoadQueue.scala 163:19:@14027.4]
  wire  storeAddrNotKnownFlags_9_10; // @[LoadQueue.scala 163:19:@14029.4]
  wire  storeAddrNotKnownFlags_9_11; // @[LoadQueue.scala 163:19:@14031.4]
  wire  storeAddrNotKnownFlags_9_12; // @[LoadQueue.scala 163:19:@14033.4]
  wire  storeAddrNotKnownFlags_9_13; // @[LoadQueue.scala 163:19:@14035.4]
  wire  storeAddrNotKnownFlags_9_14; // @[LoadQueue.scala 163:19:@14037.4]
  wire  storeAddrNotKnownFlags_9_15; // @[LoadQueue.scala 163:19:@14039.4]
  wire  storeAddrNotKnownFlags_10_0; // @[LoadQueue.scala 163:19:@14057.4]
  wire  storeAddrNotKnownFlags_10_1; // @[LoadQueue.scala 163:19:@14059.4]
  wire  storeAddrNotKnownFlags_10_2; // @[LoadQueue.scala 163:19:@14061.4]
  wire  storeAddrNotKnownFlags_10_3; // @[LoadQueue.scala 163:19:@14063.4]
  wire  storeAddrNotKnownFlags_10_4; // @[LoadQueue.scala 163:19:@14065.4]
  wire  storeAddrNotKnownFlags_10_5; // @[LoadQueue.scala 163:19:@14067.4]
  wire  storeAddrNotKnownFlags_10_6; // @[LoadQueue.scala 163:19:@14069.4]
  wire  storeAddrNotKnownFlags_10_7; // @[LoadQueue.scala 163:19:@14071.4]
  wire  storeAddrNotKnownFlags_10_8; // @[LoadQueue.scala 163:19:@14073.4]
  wire  storeAddrNotKnownFlags_10_9; // @[LoadQueue.scala 163:19:@14075.4]
  wire  storeAddrNotKnownFlags_10_10; // @[LoadQueue.scala 163:19:@14077.4]
  wire  storeAddrNotKnownFlags_10_11; // @[LoadQueue.scala 163:19:@14079.4]
  wire  storeAddrNotKnownFlags_10_12; // @[LoadQueue.scala 163:19:@14081.4]
  wire  storeAddrNotKnownFlags_10_13; // @[LoadQueue.scala 163:19:@14083.4]
  wire  storeAddrNotKnownFlags_10_14; // @[LoadQueue.scala 163:19:@14085.4]
  wire  storeAddrNotKnownFlags_10_15; // @[LoadQueue.scala 163:19:@14087.4]
  wire  storeAddrNotKnownFlags_11_0; // @[LoadQueue.scala 163:19:@14105.4]
  wire  storeAddrNotKnownFlags_11_1; // @[LoadQueue.scala 163:19:@14107.4]
  wire  storeAddrNotKnownFlags_11_2; // @[LoadQueue.scala 163:19:@14109.4]
  wire  storeAddrNotKnownFlags_11_3; // @[LoadQueue.scala 163:19:@14111.4]
  wire  storeAddrNotKnownFlags_11_4; // @[LoadQueue.scala 163:19:@14113.4]
  wire  storeAddrNotKnownFlags_11_5; // @[LoadQueue.scala 163:19:@14115.4]
  wire  storeAddrNotKnownFlags_11_6; // @[LoadQueue.scala 163:19:@14117.4]
  wire  storeAddrNotKnownFlags_11_7; // @[LoadQueue.scala 163:19:@14119.4]
  wire  storeAddrNotKnownFlags_11_8; // @[LoadQueue.scala 163:19:@14121.4]
  wire  storeAddrNotKnownFlags_11_9; // @[LoadQueue.scala 163:19:@14123.4]
  wire  storeAddrNotKnownFlags_11_10; // @[LoadQueue.scala 163:19:@14125.4]
  wire  storeAddrNotKnownFlags_11_11; // @[LoadQueue.scala 163:19:@14127.4]
  wire  storeAddrNotKnownFlags_11_12; // @[LoadQueue.scala 163:19:@14129.4]
  wire  storeAddrNotKnownFlags_11_13; // @[LoadQueue.scala 163:19:@14131.4]
  wire  storeAddrNotKnownFlags_11_14; // @[LoadQueue.scala 163:19:@14133.4]
  wire  storeAddrNotKnownFlags_11_15; // @[LoadQueue.scala 163:19:@14135.4]
  wire  storeAddrNotKnownFlags_12_0; // @[LoadQueue.scala 163:19:@14153.4]
  wire  storeAddrNotKnownFlags_12_1; // @[LoadQueue.scala 163:19:@14155.4]
  wire  storeAddrNotKnownFlags_12_2; // @[LoadQueue.scala 163:19:@14157.4]
  wire  storeAddrNotKnownFlags_12_3; // @[LoadQueue.scala 163:19:@14159.4]
  wire  storeAddrNotKnownFlags_12_4; // @[LoadQueue.scala 163:19:@14161.4]
  wire  storeAddrNotKnownFlags_12_5; // @[LoadQueue.scala 163:19:@14163.4]
  wire  storeAddrNotKnownFlags_12_6; // @[LoadQueue.scala 163:19:@14165.4]
  wire  storeAddrNotKnownFlags_12_7; // @[LoadQueue.scala 163:19:@14167.4]
  wire  storeAddrNotKnownFlags_12_8; // @[LoadQueue.scala 163:19:@14169.4]
  wire  storeAddrNotKnownFlags_12_9; // @[LoadQueue.scala 163:19:@14171.4]
  wire  storeAddrNotKnownFlags_12_10; // @[LoadQueue.scala 163:19:@14173.4]
  wire  storeAddrNotKnownFlags_12_11; // @[LoadQueue.scala 163:19:@14175.4]
  wire  storeAddrNotKnownFlags_12_12; // @[LoadQueue.scala 163:19:@14177.4]
  wire  storeAddrNotKnownFlags_12_13; // @[LoadQueue.scala 163:19:@14179.4]
  wire  storeAddrNotKnownFlags_12_14; // @[LoadQueue.scala 163:19:@14181.4]
  wire  storeAddrNotKnownFlags_12_15; // @[LoadQueue.scala 163:19:@14183.4]
  wire  storeAddrNotKnownFlags_13_0; // @[LoadQueue.scala 163:19:@14201.4]
  wire  storeAddrNotKnownFlags_13_1; // @[LoadQueue.scala 163:19:@14203.4]
  wire  storeAddrNotKnownFlags_13_2; // @[LoadQueue.scala 163:19:@14205.4]
  wire  storeAddrNotKnownFlags_13_3; // @[LoadQueue.scala 163:19:@14207.4]
  wire  storeAddrNotKnownFlags_13_4; // @[LoadQueue.scala 163:19:@14209.4]
  wire  storeAddrNotKnownFlags_13_5; // @[LoadQueue.scala 163:19:@14211.4]
  wire  storeAddrNotKnownFlags_13_6; // @[LoadQueue.scala 163:19:@14213.4]
  wire  storeAddrNotKnownFlags_13_7; // @[LoadQueue.scala 163:19:@14215.4]
  wire  storeAddrNotKnownFlags_13_8; // @[LoadQueue.scala 163:19:@14217.4]
  wire  storeAddrNotKnownFlags_13_9; // @[LoadQueue.scala 163:19:@14219.4]
  wire  storeAddrNotKnownFlags_13_10; // @[LoadQueue.scala 163:19:@14221.4]
  wire  storeAddrNotKnownFlags_13_11; // @[LoadQueue.scala 163:19:@14223.4]
  wire  storeAddrNotKnownFlags_13_12; // @[LoadQueue.scala 163:19:@14225.4]
  wire  storeAddrNotKnownFlags_13_13; // @[LoadQueue.scala 163:19:@14227.4]
  wire  storeAddrNotKnownFlags_13_14; // @[LoadQueue.scala 163:19:@14229.4]
  wire  storeAddrNotKnownFlags_13_15; // @[LoadQueue.scala 163:19:@14231.4]
  wire  storeAddrNotKnownFlags_14_0; // @[LoadQueue.scala 163:19:@14249.4]
  wire  storeAddrNotKnownFlags_14_1; // @[LoadQueue.scala 163:19:@14251.4]
  wire  storeAddrNotKnownFlags_14_2; // @[LoadQueue.scala 163:19:@14253.4]
  wire  storeAddrNotKnownFlags_14_3; // @[LoadQueue.scala 163:19:@14255.4]
  wire  storeAddrNotKnownFlags_14_4; // @[LoadQueue.scala 163:19:@14257.4]
  wire  storeAddrNotKnownFlags_14_5; // @[LoadQueue.scala 163:19:@14259.4]
  wire  storeAddrNotKnownFlags_14_6; // @[LoadQueue.scala 163:19:@14261.4]
  wire  storeAddrNotKnownFlags_14_7; // @[LoadQueue.scala 163:19:@14263.4]
  wire  storeAddrNotKnownFlags_14_8; // @[LoadQueue.scala 163:19:@14265.4]
  wire  storeAddrNotKnownFlags_14_9; // @[LoadQueue.scala 163:19:@14267.4]
  wire  storeAddrNotKnownFlags_14_10; // @[LoadQueue.scala 163:19:@14269.4]
  wire  storeAddrNotKnownFlags_14_11; // @[LoadQueue.scala 163:19:@14271.4]
  wire  storeAddrNotKnownFlags_14_12; // @[LoadQueue.scala 163:19:@14273.4]
  wire  storeAddrNotKnownFlags_14_13; // @[LoadQueue.scala 163:19:@14275.4]
  wire  storeAddrNotKnownFlags_14_14; // @[LoadQueue.scala 163:19:@14277.4]
  wire  storeAddrNotKnownFlags_14_15; // @[LoadQueue.scala 163:19:@14279.4]
  wire  storeAddrNotKnownFlags_15_0; // @[LoadQueue.scala 163:19:@14297.4]
  wire  storeAddrNotKnownFlags_15_1; // @[LoadQueue.scala 163:19:@14299.4]
  wire  storeAddrNotKnownFlags_15_2; // @[LoadQueue.scala 163:19:@14301.4]
  wire  storeAddrNotKnownFlags_15_3; // @[LoadQueue.scala 163:19:@14303.4]
  wire  storeAddrNotKnownFlags_15_4; // @[LoadQueue.scala 163:19:@14305.4]
  wire  storeAddrNotKnownFlags_15_5; // @[LoadQueue.scala 163:19:@14307.4]
  wire  storeAddrNotKnownFlags_15_6; // @[LoadQueue.scala 163:19:@14309.4]
  wire  storeAddrNotKnownFlags_15_7; // @[LoadQueue.scala 163:19:@14311.4]
  wire  storeAddrNotKnownFlags_15_8; // @[LoadQueue.scala 163:19:@14313.4]
  wire  storeAddrNotKnownFlags_15_9; // @[LoadQueue.scala 163:19:@14315.4]
  wire  storeAddrNotKnownFlags_15_10; // @[LoadQueue.scala 163:19:@14317.4]
  wire  storeAddrNotKnownFlags_15_11; // @[LoadQueue.scala 163:19:@14319.4]
  wire  storeAddrNotKnownFlags_15_12; // @[LoadQueue.scala 163:19:@14321.4]
  wire  storeAddrNotKnownFlags_15_13; // @[LoadQueue.scala 163:19:@14323.4]
  wire  storeAddrNotKnownFlags_15_14; // @[LoadQueue.scala 163:19:@14325.4]
  wire  storeAddrNotKnownFlags_15_15; // @[LoadQueue.scala 163:19:@14327.4]
  wire [7:0] _T_18002; // @[Mux.scala 19:72:@14658.4]
  wire [7:0] _T_18009; // @[Mux.scala 19:72:@14665.4]
  wire [15:0] _T_18010; // @[Mux.scala 19:72:@14666.4]
  wire [15:0] _T_18012; // @[Mux.scala 19:72:@14667.4]
  wire [7:0] _T_18019; // @[Mux.scala 19:72:@14674.4]
  wire [7:0] _T_18026; // @[Mux.scala 19:72:@14681.4]
  wire [15:0] _T_18027; // @[Mux.scala 19:72:@14682.4]
  wire [15:0] _T_18029; // @[Mux.scala 19:72:@14683.4]
  wire [7:0] _T_18036; // @[Mux.scala 19:72:@14690.4]
  wire [7:0] _T_18043; // @[Mux.scala 19:72:@14697.4]
  wire [15:0] _T_18044; // @[Mux.scala 19:72:@14698.4]
  wire [15:0] _T_18046; // @[Mux.scala 19:72:@14699.4]
  wire [7:0] _T_18053; // @[Mux.scala 19:72:@14706.4]
  wire [7:0] _T_18060; // @[Mux.scala 19:72:@14713.4]
  wire [15:0] _T_18061; // @[Mux.scala 19:72:@14714.4]
  wire [15:0] _T_18063; // @[Mux.scala 19:72:@14715.4]
  wire [7:0] _T_18070; // @[Mux.scala 19:72:@14722.4]
  wire [7:0] _T_18077; // @[Mux.scala 19:72:@14729.4]
  wire [15:0] _T_18078; // @[Mux.scala 19:72:@14730.4]
  wire [15:0] _T_18080; // @[Mux.scala 19:72:@14731.4]
  wire [7:0] _T_18087; // @[Mux.scala 19:72:@14738.4]
  wire [7:0] _T_18094; // @[Mux.scala 19:72:@14745.4]
  wire [15:0] _T_18095; // @[Mux.scala 19:72:@14746.4]
  wire [15:0] _T_18097; // @[Mux.scala 19:72:@14747.4]
  wire [7:0] _T_18104; // @[Mux.scala 19:72:@14754.4]
  wire [7:0] _T_18111; // @[Mux.scala 19:72:@14761.4]
  wire [15:0] _T_18112; // @[Mux.scala 19:72:@14762.4]
  wire [15:0] _T_18114; // @[Mux.scala 19:72:@14763.4]
  wire [7:0] _T_18121; // @[Mux.scala 19:72:@14770.4]
  wire [7:0] _T_18128; // @[Mux.scala 19:72:@14777.4]
  wire [15:0] _T_18129; // @[Mux.scala 19:72:@14778.4]
  wire [15:0] _T_18131; // @[Mux.scala 19:72:@14779.4]
  wire [15:0] _T_18146; // @[Mux.scala 19:72:@14794.4]
  wire [15:0] _T_18148; // @[Mux.scala 19:72:@14795.4]
  wire [15:0] _T_18163; // @[Mux.scala 19:72:@14810.4]
  wire [15:0] _T_18165; // @[Mux.scala 19:72:@14811.4]
  wire [15:0] _T_18180; // @[Mux.scala 19:72:@14826.4]
  wire [15:0] _T_18182; // @[Mux.scala 19:72:@14827.4]
  wire [15:0] _T_18197; // @[Mux.scala 19:72:@14842.4]
  wire [15:0] _T_18199; // @[Mux.scala 19:72:@14843.4]
  wire [15:0] _T_18214; // @[Mux.scala 19:72:@14858.4]
  wire [15:0] _T_18216; // @[Mux.scala 19:72:@14859.4]
  wire [15:0] _T_18231; // @[Mux.scala 19:72:@14874.4]
  wire [15:0] _T_18233; // @[Mux.scala 19:72:@14875.4]
  wire [15:0] _T_18248; // @[Mux.scala 19:72:@14890.4]
  wire [15:0] _T_18250; // @[Mux.scala 19:72:@14891.4]
  wire [15:0] _T_18265; // @[Mux.scala 19:72:@14906.4]
  wire [15:0] _T_18267; // @[Mux.scala 19:72:@14907.4]
  wire [15:0] _T_18268; // @[Mux.scala 19:72:@14908.4]
  wire [15:0] _T_18269; // @[Mux.scala 19:72:@14909.4]
  wire [15:0] _T_18270; // @[Mux.scala 19:72:@14910.4]
  wire [15:0] _T_18271; // @[Mux.scala 19:72:@14911.4]
  wire [15:0] _T_18272; // @[Mux.scala 19:72:@14912.4]
  wire [15:0] _T_18273; // @[Mux.scala 19:72:@14913.4]
  wire [15:0] _T_18274; // @[Mux.scala 19:72:@14914.4]
  wire [15:0] _T_18275; // @[Mux.scala 19:72:@14915.4]
  wire [15:0] _T_18276; // @[Mux.scala 19:72:@14916.4]
  wire [15:0] _T_18277; // @[Mux.scala 19:72:@14917.4]
  wire [15:0] _T_18278; // @[Mux.scala 19:72:@14918.4]
  wire [15:0] _T_18279; // @[Mux.scala 19:72:@14919.4]
  wire [15:0] _T_18280; // @[Mux.scala 19:72:@14920.4]
  wire [15:0] _T_18281; // @[Mux.scala 19:72:@14921.4]
  wire [15:0] _T_18282; // @[Mux.scala 19:72:@14922.4]
  wire [7:0] _T_18860; // @[Mux.scala 19:72:@15272.4]
  wire [7:0] _T_18867; // @[Mux.scala 19:72:@15279.4]
  wire [15:0] _T_18868; // @[Mux.scala 19:72:@15280.4]
  wire [15:0] _T_18870; // @[Mux.scala 19:72:@15281.4]
  wire [7:0] _T_18877; // @[Mux.scala 19:72:@15288.4]
  wire [7:0] _T_18884; // @[Mux.scala 19:72:@15295.4]
  wire [15:0] _T_18885; // @[Mux.scala 19:72:@15296.4]
  wire [15:0] _T_18887; // @[Mux.scala 19:72:@15297.4]
  wire [7:0] _T_18894; // @[Mux.scala 19:72:@15304.4]
  wire [7:0] _T_18901; // @[Mux.scala 19:72:@15311.4]
  wire [15:0] _T_18902; // @[Mux.scala 19:72:@15312.4]
  wire [15:0] _T_18904; // @[Mux.scala 19:72:@15313.4]
  wire [7:0] _T_18911; // @[Mux.scala 19:72:@15320.4]
  wire [7:0] _T_18918; // @[Mux.scala 19:72:@15327.4]
  wire [15:0] _T_18919; // @[Mux.scala 19:72:@15328.4]
  wire [15:0] _T_18921; // @[Mux.scala 19:72:@15329.4]
  wire [7:0] _T_18928; // @[Mux.scala 19:72:@15336.4]
  wire [7:0] _T_18935; // @[Mux.scala 19:72:@15343.4]
  wire [15:0] _T_18936; // @[Mux.scala 19:72:@15344.4]
  wire [15:0] _T_18938; // @[Mux.scala 19:72:@15345.4]
  wire [7:0] _T_18945; // @[Mux.scala 19:72:@15352.4]
  wire [7:0] _T_18952; // @[Mux.scala 19:72:@15359.4]
  wire [15:0] _T_18953; // @[Mux.scala 19:72:@15360.4]
  wire [15:0] _T_18955; // @[Mux.scala 19:72:@15361.4]
  wire [7:0] _T_18962; // @[Mux.scala 19:72:@15368.4]
  wire [7:0] _T_18969; // @[Mux.scala 19:72:@15375.4]
  wire [15:0] _T_18970; // @[Mux.scala 19:72:@15376.4]
  wire [15:0] _T_18972; // @[Mux.scala 19:72:@15377.4]
  wire [7:0] _T_18979; // @[Mux.scala 19:72:@15384.4]
  wire [7:0] _T_18986; // @[Mux.scala 19:72:@15391.4]
  wire [15:0] _T_18987; // @[Mux.scala 19:72:@15392.4]
  wire [15:0] _T_18989; // @[Mux.scala 19:72:@15393.4]
  wire [15:0] _T_19004; // @[Mux.scala 19:72:@15408.4]
  wire [15:0] _T_19006; // @[Mux.scala 19:72:@15409.4]
  wire [15:0] _T_19021; // @[Mux.scala 19:72:@15424.4]
  wire [15:0] _T_19023; // @[Mux.scala 19:72:@15425.4]
  wire [15:0] _T_19038; // @[Mux.scala 19:72:@15440.4]
  wire [15:0] _T_19040; // @[Mux.scala 19:72:@15441.4]
  wire [15:0] _T_19055; // @[Mux.scala 19:72:@15456.4]
  wire [15:0] _T_19057; // @[Mux.scala 19:72:@15457.4]
  wire [15:0] _T_19072; // @[Mux.scala 19:72:@15472.4]
  wire [15:0] _T_19074; // @[Mux.scala 19:72:@15473.4]
  wire [15:0] _T_19089; // @[Mux.scala 19:72:@15488.4]
  wire [15:0] _T_19091; // @[Mux.scala 19:72:@15489.4]
  wire [15:0] _T_19106; // @[Mux.scala 19:72:@15504.4]
  wire [15:0] _T_19108; // @[Mux.scala 19:72:@15505.4]
  wire [15:0] _T_19123; // @[Mux.scala 19:72:@15520.4]
  wire [15:0] _T_19125; // @[Mux.scala 19:72:@15521.4]
  wire [15:0] _T_19126; // @[Mux.scala 19:72:@15522.4]
  wire [15:0] _T_19127; // @[Mux.scala 19:72:@15523.4]
  wire [15:0] _T_19128; // @[Mux.scala 19:72:@15524.4]
  wire [15:0] _T_19129; // @[Mux.scala 19:72:@15525.4]
  wire [15:0] _T_19130; // @[Mux.scala 19:72:@15526.4]
  wire [15:0] _T_19131; // @[Mux.scala 19:72:@15527.4]
  wire [15:0] _T_19132; // @[Mux.scala 19:72:@15528.4]
  wire [15:0] _T_19133; // @[Mux.scala 19:72:@15529.4]
  wire [15:0] _T_19134; // @[Mux.scala 19:72:@15530.4]
  wire [15:0] _T_19135; // @[Mux.scala 19:72:@15531.4]
  wire [15:0] _T_19136; // @[Mux.scala 19:72:@15532.4]
  wire [15:0] _T_19137; // @[Mux.scala 19:72:@15533.4]
  wire [15:0] _T_19138; // @[Mux.scala 19:72:@15534.4]
  wire [15:0] _T_19139; // @[Mux.scala 19:72:@15535.4]
  wire [15:0] _T_19140; // @[Mux.scala 19:72:@15536.4]
  wire [7:0] _T_19718; // @[Mux.scala 19:72:@15886.4]
  wire [7:0] _T_19725; // @[Mux.scala 19:72:@15893.4]
  wire [15:0] _T_19726; // @[Mux.scala 19:72:@15894.4]
  wire [15:0] _T_19728; // @[Mux.scala 19:72:@15895.4]
  wire [7:0] _T_19735; // @[Mux.scala 19:72:@15902.4]
  wire [7:0] _T_19742; // @[Mux.scala 19:72:@15909.4]
  wire [15:0] _T_19743; // @[Mux.scala 19:72:@15910.4]
  wire [15:0] _T_19745; // @[Mux.scala 19:72:@15911.4]
  wire [7:0] _T_19752; // @[Mux.scala 19:72:@15918.4]
  wire [7:0] _T_19759; // @[Mux.scala 19:72:@15925.4]
  wire [15:0] _T_19760; // @[Mux.scala 19:72:@15926.4]
  wire [15:0] _T_19762; // @[Mux.scala 19:72:@15927.4]
  wire [7:0] _T_19769; // @[Mux.scala 19:72:@15934.4]
  wire [7:0] _T_19776; // @[Mux.scala 19:72:@15941.4]
  wire [15:0] _T_19777; // @[Mux.scala 19:72:@15942.4]
  wire [15:0] _T_19779; // @[Mux.scala 19:72:@15943.4]
  wire [7:0] _T_19786; // @[Mux.scala 19:72:@15950.4]
  wire [7:0] _T_19793; // @[Mux.scala 19:72:@15957.4]
  wire [15:0] _T_19794; // @[Mux.scala 19:72:@15958.4]
  wire [15:0] _T_19796; // @[Mux.scala 19:72:@15959.4]
  wire [7:0] _T_19803; // @[Mux.scala 19:72:@15966.4]
  wire [7:0] _T_19810; // @[Mux.scala 19:72:@15973.4]
  wire [15:0] _T_19811; // @[Mux.scala 19:72:@15974.4]
  wire [15:0] _T_19813; // @[Mux.scala 19:72:@15975.4]
  wire [7:0] _T_19820; // @[Mux.scala 19:72:@15982.4]
  wire [7:0] _T_19827; // @[Mux.scala 19:72:@15989.4]
  wire [15:0] _T_19828; // @[Mux.scala 19:72:@15990.4]
  wire [15:0] _T_19830; // @[Mux.scala 19:72:@15991.4]
  wire [7:0] _T_19837; // @[Mux.scala 19:72:@15998.4]
  wire [7:0] _T_19844; // @[Mux.scala 19:72:@16005.4]
  wire [15:0] _T_19845; // @[Mux.scala 19:72:@16006.4]
  wire [15:0] _T_19847; // @[Mux.scala 19:72:@16007.4]
  wire [15:0] _T_19862; // @[Mux.scala 19:72:@16022.4]
  wire [15:0] _T_19864; // @[Mux.scala 19:72:@16023.4]
  wire [15:0] _T_19879; // @[Mux.scala 19:72:@16038.4]
  wire [15:0] _T_19881; // @[Mux.scala 19:72:@16039.4]
  wire [15:0] _T_19896; // @[Mux.scala 19:72:@16054.4]
  wire [15:0] _T_19898; // @[Mux.scala 19:72:@16055.4]
  wire [15:0] _T_19913; // @[Mux.scala 19:72:@16070.4]
  wire [15:0] _T_19915; // @[Mux.scala 19:72:@16071.4]
  wire [15:0] _T_19930; // @[Mux.scala 19:72:@16086.4]
  wire [15:0] _T_19932; // @[Mux.scala 19:72:@16087.4]
  wire [15:0] _T_19947; // @[Mux.scala 19:72:@16102.4]
  wire [15:0] _T_19949; // @[Mux.scala 19:72:@16103.4]
  wire [15:0] _T_19964; // @[Mux.scala 19:72:@16118.4]
  wire [15:0] _T_19966; // @[Mux.scala 19:72:@16119.4]
  wire [15:0] _T_19981; // @[Mux.scala 19:72:@16134.4]
  wire [15:0] _T_19983; // @[Mux.scala 19:72:@16135.4]
  wire [15:0] _T_19984; // @[Mux.scala 19:72:@16136.4]
  wire [15:0] _T_19985; // @[Mux.scala 19:72:@16137.4]
  wire [15:0] _T_19986; // @[Mux.scala 19:72:@16138.4]
  wire [15:0] _T_19987; // @[Mux.scala 19:72:@16139.4]
  wire [15:0] _T_19988; // @[Mux.scala 19:72:@16140.4]
  wire [15:0] _T_19989; // @[Mux.scala 19:72:@16141.4]
  wire [15:0] _T_19990; // @[Mux.scala 19:72:@16142.4]
  wire [15:0] _T_19991; // @[Mux.scala 19:72:@16143.4]
  wire [15:0] _T_19992; // @[Mux.scala 19:72:@16144.4]
  wire [15:0] _T_19993; // @[Mux.scala 19:72:@16145.4]
  wire [15:0] _T_19994; // @[Mux.scala 19:72:@16146.4]
  wire [15:0] _T_19995; // @[Mux.scala 19:72:@16147.4]
  wire [15:0] _T_19996; // @[Mux.scala 19:72:@16148.4]
  wire [15:0] _T_19997; // @[Mux.scala 19:72:@16149.4]
  wire [15:0] _T_19998; // @[Mux.scala 19:72:@16150.4]
  wire [7:0] _T_20576; // @[Mux.scala 19:72:@16500.4]
  wire [7:0] _T_20583; // @[Mux.scala 19:72:@16507.4]
  wire [15:0] _T_20584; // @[Mux.scala 19:72:@16508.4]
  wire [15:0] _T_20586; // @[Mux.scala 19:72:@16509.4]
  wire [7:0] _T_20593; // @[Mux.scala 19:72:@16516.4]
  wire [7:0] _T_20600; // @[Mux.scala 19:72:@16523.4]
  wire [15:0] _T_20601; // @[Mux.scala 19:72:@16524.4]
  wire [15:0] _T_20603; // @[Mux.scala 19:72:@16525.4]
  wire [7:0] _T_20610; // @[Mux.scala 19:72:@16532.4]
  wire [7:0] _T_20617; // @[Mux.scala 19:72:@16539.4]
  wire [15:0] _T_20618; // @[Mux.scala 19:72:@16540.4]
  wire [15:0] _T_20620; // @[Mux.scala 19:72:@16541.4]
  wire [7:0] _T_20627; // @[Mux.scala 19:72:@16548.4]
  wire [7:0] _T_20634; // @[Mux.scala 19:72:@16555.4]
  wire [15:0] _T_20635; // @[Mux.scala 19:72:@16556.4]
  wire [15:0] _T_20637; // @[Mux.scala 19:72:@16557.4]
  wire [7:0] _T_20644; // @[Mux.scala 19:72:@16564.4]
  wire [7:0] _T_20651; // @[Mux.scala 19:72:@16571.4]
  wire [15:0] _T_20652; // @[Mux.scala 19:72:@16572.4]
  wire [15:0] _T_20654; // @[Mux.scala 19:72:@16573.4]
  wire [7:0] _T_20661; // @[Mux.scala 19:72:@16580.4]
  wire [7:0] _T_20668; // @[Mux.scala 19:72:@16587.4]
  wire [15:0] _T_20669; // @[Mux.scala 19:72:@16588.4]
  wire [15:0] _T_20671; // @[Mux.scala 19:72:@16589.4]
  wire [7:0] _T_20678; // @[Mux.scala 19:72:@16596.4]
  wire [7:0] _T_20685; // @[Mux.scala 19:72:@16603.4]
  wire [15:0] _T_20686; // @[Mux.scala 19:72:@16604.4]
  wire [15:0] _T_20688; // @[Mux.scala 19:72:@16605.4]
  wire [7:0] _T_20695; // @[Mux.scala 19:72:@16612.4]
  wire [7:0] _T_20702; // @[Mux.scala 19:72:@16619.4]
  wire [15:0] _T_20703; // @[Mux.scala 19:72:@16620.4]
  wire [15:0] _T_20705; // @[Mux.scala 19:72:@16621.4]
  wire [15:0] _T_20720; // @[Mux.scala 19:72:@16636.4]
  wire [15:0] _T_20722; // @[Mux.scala 19:72:@16637.4]
  wire [15:0] _T_20737; // @[Mux.scala 19:72:@16652.4]
  wire [15:0] _T_20739; // @[Mux.scala 19:72:@16653.4]
  wire [15:0] _T_20754; // @[Mux.scala 19:72:@16668.4]
  wire [15:0] _T_20756; // @[Mux.scala 19:72:@16669.4]
  wire [15:0] _T_20771; // @[Mux.scala 19:72:@16684.4]
  wire [15:0] _T_20773; // @[Mux.scala 19:72:@16685.4]
  wire [15:0] _T_20788; // @[Mux.scala 19:72:@16700.4]
  wire [15:0] _T_20790; // @[Mux.scala 19:72:@16701.4]
  wire [15:0] _T_20805; // @[Mux.scala 19:72:@16716.4]
  wire [15:0] _T_20807; // @[Mux.scala 19:72:@16717.4]
  wire [15:0] _T_20822; // @[Mux.scala 19:72:@16732.4]
  wire [15:0] _T_20824; // @[Mux.scala 19:72:@16733.4]
  wire [15:0] _T_20839; // @[Mux.scala 19:72:@16748.4]
  wire [15:0] _T_20841; // @[Mux.scala 19:72:@16749.4]
  wire [15:0] _T_20842; // @[Mux.scala 19:72:@16750.4]
  wire [15:0] _T_20843; // @[Mux.scala 19:72:@16751.4]
  wire [15:0] _T_20844; // @[Mux.scala 19:72:@16752.4]
  wire [15:0] _T_20845; // @[Mux.scala 19:72:@16753.4]
  wire [15:0] _T_20846; // @[Mux.scala 19:72:@16754.4]
  wire [15:0] _T_20847; // @[Mux.scala 19:72:@16755.4]
  wire [15:0] _T_20848; // @[Mux.scala 19:72:@16756.4]
  wire [15:0] _T_20849; // @[Mux.scala 19:72:@16757.4]
  wire [15:0] _T_20850; // @[Mux.scala 19:72:@16758.4]
  wire [15:0] _T_20851; // @[Mux.scala 19:72:@16759.4]
  wire [15:0] _T_20852; // @[Mux.scala 19:72:@16760.4]
  wire [15:0] _T_20853; // @[Mux.scala 19:72:@16761.4]
  wire [15:0] _T_20854; // @[Mux.scala 19:72:@16762.4]
  wire [15:0] _T_20855; // @[Mux.scala 19:72:@16763.4]
  wire [15:0] _T_20856; // @[Mux.scala 19:72:@16764.4]
  wire [7:0] _T_21434; // @[Mux.scala 19:72:@17114.4]
  wire [7:0] _T_21441; // @[Mux.scala 19:72:@17121.4]
  wire [15:0] _T_21442; // @[Mux.scala 19:72:@17122.4]
  wire [15:0] _T_21444; // @[Mux.scala 19:72:@17123.4]
  wire [7:0] _T_21451; // @[Mux.scala 19:72:@17130.4]
  wire [7:0] _T_21458; // @[Mux.scala 19:72:@17137.4]
  wire [15:0] _T_21459; // @[Mux.scala 19:72:@17138.4]
  wire [15:0] _T_21461; // @[Mux.scala 19:72:@17139.4]
  wire [7:0] _T_21468; // @[Mux.scala 19:72:@17146.4]
  wire [7:0] _T_21475; // @[Mux.scala 19:72:@17153.4]
  wire [15:0] _T_21476; // @[Mux.scala 19:72:@17154.4]
  wire [15:0] _T_21478; // @[Mux.scala 19:72:@17155.4]
  wire [7:0] _T_21485; // @[Mux.scala 19:72:@17162.4]
  wire [7:0] _T_21492; // @[Mux.scala 19:72:@17169.4]
  wire [15:0] _T_21493; // @[Mux.scala 19:72:@17170.4]
  wire [15:0] _T_21495; // @[Mux.scala 19:72:@17171.4]
  wire [7:0] _T_21502; // @[Mux.scala 19:72:@17178.4]
  wire [7:0] _T_21509; // @[Mux.scala 19:72:@17185.4]
  wire [15:0] _T_21510; // @[Mux.scala 19:72:@17186.4]
  wire [15:0] _T_21512; // @[Mux.scala 19:72:@17187.4]
  wire [7:0] _T_21519; // @[Mux.scala 19:72:@17194.4]
  wire [7:0] _T_21526; // @[Mux.scala 19:72:@17201.4]
  wire [15:0] _T_21527; // @[Mux.scala 19:72:@17202.4]
  wire [15:0] _T_21529; // @[Mux.scala 19:72:@17203.4]
  wire [7:0] _T_21536; // @[Mux.scala 19:72:@17210.4]
  wire [7:0] _T_21543; // @[Mux.scala 19:72:@17217.4]
  wire [15:0] _T_21544; // @[Mux.scala 19:72:@17218.4]
  wire [15:0] _T_21546; // @[Mux.scala 19:72:@17219.4]
  wire [7:0] _T_21553; // @[Mux.scala 19:72:@17226.4]
  wire [7:0] _T_21560; // @[Mux.scala 19:72:@17233.4]
  wire [15:0] _T_21561; // @[Mux.scala 19:72:@17234.4]
  wire [15:0] _T_21563; // @[Mux.scala 19:72:@17235.4]
  wire [15:0] _T_21578; // @[Mux.scala 19:72:@17250.4]
  wire [15:0] _T_21580; // @[Mux.scala 19:72:@17251.4]
  wire [15:0] _T_21595; // @[Mux.scala 19:72:@17266.4]
  wire [15:0] _T_21597; // @[Mux.scala 19:72:@17267.4]
  wire [15:0] _T_21612; // @[Mux.scala 19:72:@17282.4]
  wire [15:0] _T_21614; // @[Mux.scala 19:72:@17283.4]
  wire [15:0] _T_21629; // @[Mux.scala 19:72:@17298.4]
  wire [15:0] _T_21631; // @[Mux.scala 19:72:@17299.4]
  wire [15:0] _T_21646; // @[Mux.scala 19:72:@17314.4]
  wire [15:0] _T_21648; // @[Mux.scala 19:72:@17315.4]
  wire [15:0] _T_21663; // @[Mux.scala 19:72:@17330.4]
  wire [15:0] _T_21665; // @[Mux.scala 19:72:@17331.4]
  wire [15:0] _T_21680; // @[Mux.scala 19:72:@17346.4]
  wire [15:0] _T_21682; // @[Mux.scala 19:72:@17347.4]
  wire [15:0] _T_21697; // @[Mux.scala 19:72:@17362.4]
  wire [15:0] _T_21699; // @[Mux.scala 19:72:@17363.4]
  wire [15:0] _T_21700; // @[Mux.scala 19:72:@17364.4]
  wire [15:0] _T_21701; // @[Mux.scala 19:72:@17365.4]
  wire [15:0] _T_21702; // @[Mux.scala 19:72:@17366.4]
  wire [15:0] _T_21703; // @[Mux.scala 19:72:@17367.4]
  wire [15:0] _T_21704; // @[Mux.scala 19:72:@17368.4]
  wire [15:0] _T_21705; // @[Mux.scala 19:72:@17369.4]
  wire [15:0] _T_21706; // @[Mux.scala 19:72:@17370.4]
  wire [15:0] _T_21707; // @[Mux.scala 19:72:@17371.4]
  wire [15:0] _T_21708; // @[Mux.scala 19:72:@17372.4]
  wire [15:0] _T_21709; // @[Mux.scala 19:72:@17373.4]
  wire [15:0] _T_21710; // @[Mux.scala 19:72:@17374.4]
  wire [15:0] _T_21711; // @[Mux.scala 19:72:@17375.4]
  wire [15:0] _T_21712; // @[Mux.scala 19:72:@17376.4]
  wire [15:0] _T_21713; // @[Mux.scala 19:72:@17377.4]
  wire [15:0] _T_21714; // @[Mux.scala 19:72:@17378.4]
  wire [7:0] _T_22292; // @[Mux.scala 19:72:@17728.4]
  wire [7:0] _T_22299; // @[Mux.scala 19:72:@17735.4]
  wire [15:0] _T_22300; // @[Mux.scala 19:72:@17736.4]
  wire [15:0] _T_22302; // @[Mux.scala 19:72:@17737.4]
  wire [7:0] _T_22309; // @[Mux.scala 19:72:@17744.4]
  wire [7:0] _T_22316; // @[Mux.scala 19:72:@17751.4]
  wire [15:0] _T_22317; // @[Mux.scala 19:72:@17752.4]
  wire [15:0] _T_22319; // @[Mux.scala 19:72:@17753.4]
  wire [7:0] _T_22326; // @[Mux.scala 19:72:@17760.4]
  wire [7:0] _T_22333; // @[Mux.scala 19:72:@17767.4]
  wire [15:0] _T_22334; // @[Mux.scala 19:72:@17768.4]
  wire [15:0] _T_22336; // @[Mux.scala 19:72:@17769.4]
  wire [7:0] _T_22343; // @[Mux.scala 19:72:@17776.4]
  wire [7:0] _T_22350; // @[Mux.scala 19:72:@17783.4]
  wire [15:0] _T_22351; // @[Mux.scala 19:72:@17784.4]
  wire [15:0] _T_22353; // @[Mux.scala 19:72:@17785.4]
  wire [7:0] _T_22360; // @[Mux.scala 19:72:@17792.4]
  wire [7:0] _T_22367; // @[Mux.scala 19:72:@17799.4]
  wire [15:0] _T_22368; // @[Mux.scala 19:72:@17800.4]
  wire [15:0] _T_22370; // @[Mux.scala 19:72:@17801.4]
  wire [7:0] _T_22377; // @[Mux.scala 19:72:@17808.4]
  wire [7:0] _T_22384; // @[Mux.scala 19:72:@17815.4]
  wire [15:0] _T_22385; // @[Mux.scala 19:72:@17816.4]
  wire [15:0] _T_22387; // @[Mux.scala 19:72:@17817.4]
  wire [7:0] _T_22394; // @[Mux.scala 19:72:@17824.4]
  wire [7:0] _T_22401; // @[Mux.scala 19:72:@17831.4]
  wire [15:0] _T_22402; // @[Mux.scala 19:72:@17832.4]
  wire [15:0] _T_22404; // @[Mux.scala 19:72:@17833.4]
  wire [7:0] _T_22411; // @[Mux.scala 19:72:@17840.4]
  wire [7:0] _T_22418; // @[Mux.scala 19:72:@17847.4]
  wire [15:0] _T_22419; // @[Mux.scala 19:72:@17848.4]
  wire [15:0] _T_22421; // @[Mux.scala 19:72:@17849.4]
  wire [15:0] _T_22436; // @[Mux.scala 19:72:@17864.4]
  wire [15:0] _T_22438; // @[Mux.scala 19:72:@17865.4]
  wire [15:0] _T_22453; // @[Mux.scala 19:72:@17880.4]
  wire [15:0] _T_22455; // @[Mux.scala 19:72:@17881.4]
  wire [15:0] _T_22470; // @[Mux.scala 19:72:@17896.4]
  wire [15:0] _T_22472; // @[Mux.scala 19:72:@17897.4]
  wire [15:0] _T_22487; // @[Mux.scala 19:72:@17912.4]
  wire [15:0] _T_22489; // @[Mux.scala 19:72:@17913.4]
  wire [15:0] _T_22504; // @[Mux.scala 19:72:@17928.4]
  wire [15:0] _T_22506; // @[Mux.scala 19:72:@17929.4]
  wire [15:0] _T_22521; // @[Mux.scala 19:72:@17944.4]
  wire [15:0] _T_22523; // @[Mux.scala 19:72:@17945.4]
  wire [15:0] _T_22538; // @[Mux.scala 19:72:@17960.4]
  wire [15:0] _T_22540; // @[Mux.scala 19:72:@17961.4]
  wire [15:0] _T_22555; // @[Mux.scala 19:72:@17976.4]
  wire [15:0] _T_22557; // @[Mux.scala 19:72:@17977.4]
  wire [15:0] _T_22558; // @[Mux.scala 19:72:@17978.4]
  wire [15:0] _T_22559; // @[Mux.scala 19:72:@17979.4]
  wire [15:0] _T_22560; // @[Mux.scala 19:72:@17980.4]
  wire [15:0] _T_22561; // @[Mux.scala 19:72:@17981.4]
  wire [15:0] _T_22562; // @[Mux.scala 19:72:@17982.4]
  wire [15:0] _T_22563; // @[Mux.scala 19:72:@17983.4]
  wire [15:0] _T_22564; // @[Mux.scala 19:72:@17984.4]
  wire [15:0] _T_22565; // @[Mux.scala 19:72:@17985.4]
  wire [15:0] _T_22566; // @[Mux.scala 19:72:@17986.4]
  wire [15:0] _T_22567; // @[Mux.scala 19:72:@17987.4]
  wire [15:0] _T_22568; // @[Mux.scala 19:72:@17988.4]
  wire [15:0] _T_22569; // @[Mux.scala 19:72:@17989.4]
  wire [15:0] _T_22570; // @[Mux.scala 19:72:@17990.4]
  wire [15:0] _T_22571; // @[Mux.scala 19:72:@17991.4]
  wire [15:0] _T_22572; // @[Mux.scala 19:72:@17992.4]
  wire [7:0] _T_23150; // @[Mux.scala 19:72:@18342.4]
  wire [7:0] _T_23157; // @[Mux.scala 19:72:@18349.4]
  wire [15:0] _T_23158; // @[Mux.scala 19:72:@18350.4]
  wire [15:0] _T_23160; // @[Mux.scala 19:72:@18351.4]
  wire [7:0] _T_23167; // @[Mux.scala 19:72:@18358.4]
  wire [7:0] _T_23174; // @[Mux.scala 19:72:@18365.4]
  wire [15:0] _T_23175; // @[Mux.scala 19:72:@18366.4]
  wire [15:0] _T_23177; // @[Mux.scala 19:72:@18367.4]
  wire [7:0] _T_23184; // @[Mux.scala 19:72:@18374.4]
  wire [7:0] _T_23191; // @[Mux.scala 19:72:@18381.4]
  wire [15:0] _T_23192; // @[Mux.scala 19:72:@18382.4]
  wire [15:0] _T_23194; // @[Mux.scala 19:72:@18383.4]
  wire [7:0] _T_23201; // @[Mux.scala 19:72:@18390.4]
  wire [7:0] _T_23208; // @[Mux.scala 19:72:@18397.4]
  wire [15:0] _T_23209; // @[Mux.scala 19:72:@18398.4]
  wire [15:0] _T_23211; // @[Mux.scala 19:72:@18399.4]
  wire [7:0] _T_23218; // @[Mux.scala 19:72:@18406.4]
  wire [7:0] _T_23225; // @[Mux.scala 19:72:@18413.4]
  wire [15:0] _T_23226; // @[Mux.scala 19:72:@18414.4]
  wire [15:0] _T_23228; // @[Mux.scala 19:72:@18415.4]
  wire [7:0] _T_23235; // @[Mux.scala 19:72:@18422.4]
  wire [7:0] _T_23242; // @[Mux.scala 19:72:@18429.4]
  wire [15:0] _T_23243; // @[Mux.scala 19:72:@18430.4]
  wire [15:0] _T_23245; // @[Mux.scala 19:72:@18431.4]
  wire [7:0] _T_23252; // @[Mux.scala 19:72:@18438.4]
  wire [7:0] _T_23259; // @[Mux.scala 19:72:@18445.4]
  wire [15:0] _T_23260; // @[Mux.scala 19:72:@18446.4]
  wire [15:0] _T_23262; // @[Mux.scala 19:72:@18447.4]
  wire [7:0] _T_23269; // @[Mux.scala 19:72:@18454.4]
  wire [7:0] _T_23276; // @[Mux.scala 19:72:@18461.4]
  wire [15:0] _T_23277; // @[Mux.scala 19:72:@18462.4]
  wire [15:0] _T_23279; // @[Mux.scala 19:72:@18463.4]
  wire [15:0] _T_23294; // @[Mux.scala 19:72:@18478.4]
  wire [15:0] _T_23296; // @[Mux.scala 19:72:@18479.4]
  wire [15:0] _T_23311; // @[Mux.scala 19:72:@18494.4]
  wire [15:0] _T_23313; // @[Mux.scala 19:72:@18495.4]
  wire [15:0] _T_23328; // @[Mux.scala 19:72:@18510.4]
  wire [15:0] _T_23330; // @[Mux.scala 19:72:@18511.4]
  wire [15:0] _T_23345; // @[Mux.scala 19:72:@18526.4]
  wire [15:0] _T_23347; // @[Mux.scala 19:72:@18527.4]
  wire [15:0] _T_23362; // @[Mux.scala 19:72:@18542.4]
  wire [15:0] _T_23364; // @[Mux.scala 19:72:@18543.4]
  wire [15:0] _T_23379; // @[Mux.scala 19:72:@18558.4]
  wire [15:0] _T_23381; // @[Mux.scala 19:72:@18559.4]
  wire [15:0] _T_23396; // @[Mux.scala 19:72:@18574.4]
  wire [15:0] _T_23398; // @[Mux.scala 19:72:@18575.4]
  wire [15:0] _T_23413; // @[Mux.scala 19:72:@18590.4]
  wire [15:0] _T_23415; // @[Mux.scala 19:72:@18591.4]
  wire [15:0] _T_23416; // @[Mux.scala 19:72:@18592.4]
  wire [15:0] _T_23417; // @[Mux.scala 19:72:@18593.4]
  wire [15:0] _T_23418; // @[Mux.scala 19:72:@18594.4]
  wire [15:0] _T_23419; // @[Mux.scala 19:72:@18595.4]
  wire [15:0] _T_23420; // @[Mux.scala 19:72:@18596.4]
  wire [15:0] _T_23421; // @[Mux.scala 19:72:@18597.4]
  wire [15:0] _T_23422; // @[Mux.scala 19:72:@18598.4]
  wire [15:0] _T_23423; // @[Mux.scala 19:72:@18599.4]
  wire [15:0] _T_23424; // @[Mux.scala 19:72:@18600.4]
  wire [15:0] _T_23425; // @[Mux.scala 19:72:@18601.4]
  wire [15:0] _T_23426; // @[Mux.scala 19:72:@18602.4]
  wire [15:0] _T_23427; // @[Mux.scala 19:72:@18603.4]
  wire [15:0] _T_23428; // @[Mux.scala 19:72:@18604.4]
  wire [15:0] _T_23429; // @[Mux.scala 19:72:@18605.4]
  wire [15:0] _T_23430; // @[Mux.scala 19:72:@18606.4]
  wire [7:0] _T_24008; // @[Mux.scala 19:72:@18956.4]
  wire [7:0] _T_24015; // @[Mux.scala 19:72:@18963.4]
  wire [15:0] _T_24016; // @[Mux.scala 19:72:@18964.4]
  wire [15:0] _T_24018; // @[Mux.scala 19:72:@18965.4]
  wire [7:0] _T_24025; // @[Mux.scala 19:72:@18972.4]
  wire [7:0] _T_24032; // @[Mux.scala 19:72:@18979.4]
  wire [15:0] _T_24033; // @[Mux.scala 19:72:@18980.4]
  wire [15:0] _T_24035; // @[Mux.scala 19:72:@18981.4]
  wire [7:0] _T_24042; // @[Mux.scala 19:72:@18988.4]
  wire [7:0] _T_24049; // @[Mux.scala 19:72:@18995.4]
  wire [15:0] _T_24050; // @[Mux.scala 19:72:@18996.4]
  wire [15:0] _T_24052; // @[Mux.scala 19:72:@18997.4]
  wire [7:0] _T_24059; // @[Mux.scala 19:72:@19004.4]
  wire [7:0] _T_24066; // @[Mux.scala 19:72:@19011.4]
  wire [15:0] _T_24067; // @[Mux.scala 19:72:@19012.4]
  wire [15:0] _T_24069; // @[Mux.scala 19:72:@19013.4]
  wire [7:0] _T_24076; // @[Mux.scala 19:72:@19020.4]
  wire [7:0] _T_24083; // @[Mux.scala 19:72:@19027.4]
  wire [15:0] _T_24084; // @[Mux.scala 19:72:@19028.4]
  wire [15:0] _T_24086; // @[Mux.scala 19:72:@19029.4]
  wire [7:0] _T_24093; // @[Mux.scala 19:72:@19036.4]
  wire [7:0] _T_24100; // @[Mux.scala 19:72:@19043.4]
  wire [15:0] _T_24101; // @[Mux.scala 19:72:@19044.4]
  wire [15:0] _T_24103; // @[Mux.scala 19:72:@19045.4]
  wire [7:0] _T_24110; // @[Mux.scala 19:72:@19052.4]
  wire [7:0] _T_24117; // @[Mux.scala 19:72:@19059.4]
  wire [15:0] _T_24118; // @[Mux.scala 19:72:@19060.4]
  wire [15:0] _T_24120; // @[Mux.scala 19:72:@19061.4]
  wire [7:0] _T_24127; // @[Mux.scala 19:72:@19068.4]
  wire [7:0] _T_24134; // @[Mux.scala 19:72:@19075.4]
  wire [15:0] _T_24135; // @[Mux.scala 19:72:@19076.4]
  wire [15:0] _T_24137; // @[Mux.scala 19:72:@19077.4]
  wire [15:0] _T_24152; // @[Mux.scala 19:72:@19092.4]
  wire [15:0] _T_24154; // @[Mux.scala 19:72:@19093.4]
  wire [15:0] _T_24169; // @[Mux.scala 19:72:@19108.4]
  wire [15:0] _T_24171; // @[Mux.scala 19:72:@19109.4]
  wire [15:0] _T_24186; // @[Mux.scala 19:72:@19124.4]
  wire [15:0] _T_24188; // @[Mux.scala 19:72:@19125.4]
  wire [15:0] _T_24203; // @[Mux.scala 19:72:@19140.4]
  wire [15:0] _T_24205; // @[Mux.scala 19:72:@19141.4]
  wire [15:0] _T_24220; // @[Mux.scala 19:72:@19156.4]
  wire [15:0] _T_24222; // @[Mux.scala 19:72:@19157.4]
  wire [15:0] _T_24237; // @[Mux.scala 19:72:@19172.4]
  wire [15:0] _T_24239; // @[Mux.scala 19:72:@19173.4]
  wire [15:0] _T_24254; // @[Mux.scala 19:72:@19188.4]
  wire [15:0] _T_24256; // @[Mux.scala 19:72:@19189.4]
  wire [15:0] _T_24271; // @[Mux.scala 19:72:@19204.4]
  wire [15:0] _T_24273; // @[Mux.scala 19:72:@19205.4]
  wire [15:0] _T_24274; // @[Mux.scala 19:72:@19206.4]
  wire [15:0] _T_24275; // @[Mux.scala 19:72:@19207.4]
  wire [15:0] _T_24276; // @[Mux.scala 19:72:@19208.4]
  wire [15:0] _T_24277; // @[Mux.scala 19:72:@19209.4]
  wire [15:0] _T_24278; // @[Mux.scala 19:72:@19210.4]
  wire [15:0] _T_24279; // @[Mux.scala 19:72:@19211.4]
  wire [15:0] _T_24280; // @[Mux.scala 19:72:@19212.4]
  wire [15:0] _T_24281; // @[Mux.scala 19:72:@19213.4]
  wire [15:0] _T_24282; // @[Mux.scala 19:72:@19214.4]
  wire [15:0] _T_24283; // @[Mux.scala 19:72:@19215.4]
  wire [15:0] _T_24284; // @[Mux.scala 19:72:@19216.4]
  wire [15:0] _T_24285; // @[Mux.scala 19:72:@19217.4]
  wire [15:0] _T_24286; // @[Mux.scala 19:72:@19218.4]
  wire [15:0] _T_24287; // @[Mux.scala 19:72:@19219.4]
  wire [15:0] _T_24288; // @[Mux.scala 19:72:@19220.4]
  wire [7:0] _T_24866; // @[Mux.scala 19:72:@19570.4]
  wire [7:0] _T_24873; // @[Mux.scala 19:72:@19577.4]
  wire [15:0] _T_24874; // @[Mux.scala 19:72:@19578.4]
  wire [15:0] _T_24876; // @[Mux.scala 19:72:@19579.4]
  wire [7:0] _T_24883; // @[Mux.scala 19:72:@19586.4]
  wire [7:0] _T_24890; // @[Mux.scala 19:72:@19593.4]
  wire [15:0] _T_24891; // @[Mux.scala 19:72:@19594.4]
  wire [15:0] _T_24893; // @[Mux.scala 19:72:@19595.4]
  wire [7:0] _T_24900; // @[Mux.scala 19:72:@19602.4]
  wire [7:0] _T_24907; // @[Mux.scala 19:72:@19609.4]
  wire [15:0] _T_24908; // @[Mux.scala 19:72:@19610.4]
  wire [15:0] _T_24910; // @[Mux.scala 19:72:@19611.4]
  wire [7:0] _T_24917; // @[Mux.scala 19:72:@19618.4]
  wire [7:0] _T_24924; // @[Mux.scala 19:72:@19625.4]
  wire [15:0] _T_24925; // @[Mux.scala 19:72:@19626.4]
  wire [15:0] _T_24927; // @[Mux.scala 19:72:@19627.4]
  wire [7:0] _T_24934; // @[Mux.scala 19:72:@19634.4]
  wire [7:0] _T_24941; // @[Mux.scala 19:72:@19641.4]
  wire [15:0] _T_24942; // @[Mux.scala 19:72:@19642.4]
  wire [15:0] _T_24944; // @[Mux.scala 19:72:@19643.4]
  wire [7:0] _T_24951; // @[Mux.scala 19:72:@19650.4]
  wire [7:0] _T_24958; // @[Mux.scala 19:72:@19657.4]
  wire [15:0] _T_24959; // @[Mux.scala 19:72:@19658.4]
  wire [15:0] _T_24961; // @[Mux.scala 19:72:@19659.4]
  wire [7:0] _T_24968; // @[Mux.scala 19:72:@19666.4]
  wire [7:0] _T_24975; // @[Mux.scala 19:72:@19673.4]
  wire [15:0] _T_24976; // @[Mux.scala 19:72:@19674.4]
  wire [15:0] _T_24978; // @[Mux.scala 19:72:@19675.4]
  wire [7:0] _T_24985; // @[Mux.scala 19:72:@19682.4]
  wire [7:0] _T_24992; // @[Mux.scala 19:72:@19689.4]
  wire [15:0] _T_24993; // @[Mux.scala 19:72:@19690.4]
  wire [15:0] _T_24995; // @[Mux.scala 19:72:@19691.4]
  wire [15:0] _T_25010; // @[Mux.scala 19:72:@19706.4]
  wire [15:0] _T_25012; // @[Mux.scala 19:72:@19707.4]
  wire [15:0] _T_25027; // @[Mux.scala 19:72:@19722.4]
  wire [15:0] _T_25029; // @[Mux.scala 19:72:@19723.4]
  wire [15:0] _T_25044; // @[Mux.scala 19:72:@19738.4]
  wire [15:0] _T_25046; // @[Mux.scala 19:72:@19739.4]
  wire [15:0] _T_25061; // @[Mux.scala 19:72:@19754.4]
  wire [15:0] _T_25063; // @[Mux.scala 19:72:@19755.4]
  wire [15:0] _T_25078; // @[Mux.scala 19:72:@19770.4]
  wire [15:0] _T_25080; // @[Mux.scala 19:72:@19771.4]
  wire [15:0] _T_25095; // @[Mux.scala 19:72:@19786.4]
  wire [15:0] _T_25097; // @[Mux.scala 19:72:@19787.4]
  wire [15:0] _T_25112; // @[Mux.scala 19:72:@19802.4]
  wire [15:0] _T_25114; // @[Mux.scala 19:72:@19803.4]
  wire [15:0] _T_25129; // @[Mux.scala 19:72:@19818.4]
  wire [15:0] _T_25131; // @[Mux.scala 19:72:@19819.4]
  wire [15:0] _T_25132; // @[Mux.scala 19:72:@19820.4]
  wire [15:0] _T_25133; // @[Mux.scala 19:72:@19821.4]
  wire [15:0] _T_25134; // @[Mux.scala 19:72:@19822.4]
  wire [15:0] _T_25135; // @[Mux.scala 19:72:@19823.4]
  wire [15:0] _T_25136; // @[Mux.scala 19:72:@19824.4]
  wire [15:0] _T_25137; // @[Mux.scala 19:72:@19825.4]
  wire [15:0] _T_25138; // @[Mux.scala 19:72:@19826.4]
  wire [15:0] _T_25139; // @[Mux.scala 19:72:@19827.4]
  wire [15:0] _T_25140; // @[Mux.scala 19:72:@19828.4]
  wire [15:0] _T_25141; // @[Mux.scala 19:72:@19829.4]
  wire [15:0] _T_25142; // @[Mux.scala 19:72:@19830.4]
  wire [15:0] _T_25143; // @[Mux.scala 19:72:@19831.4]
  wire [15:0] _T_25144; // @[Mux.scala 19:72:@19832.4]
  wire [15:0] _T_25145; // @[Mux.scala 19:72:@19833.4]
  wire [15:0] _T_25146; // @[Mux.scala 19:72:@19834.4]
  wire [7:0] _T_25724; // @[Mux.scala 19:72:@20184.4]
  wire [7:0] _T_25731; // @[Mux.scala 19:72:@20191.4]
  wire [15:0] _T_25732; // @[Mux.scala 19:72:@20192.4]
  wire [15:0] _T_25734; // @[Mux.scala 19:72:@20193.4]
  wire [7:0] _T_25741; // @[Mux.scala 19:72:@20200.4]
  wire [7:0] _T_25748; // @[Mux.scala 19:72:@20207.4]
  wire [15:0] _T_25749; // @[Mux.scala 19:72:@20208.4]
  wire [15:0] _T_25751; // @[Mux.scala 19:72:@20209.4]
  wire [7:0] _T_25758; // @[Mux.scala 19:72:@20216.4]
  wire [7:0] _T_25765; // @[Mux.scala 19:72:@20223.4]
  wire [15:0] _T_25766; // @[Mux.scala 19:72:@20224.4]
  wire [15:0] _T_25768; // @[Mux.scala 19:72:@20225.4]
  wire [7:0] _T_25775; // @[Mux.scala 19:72:@20232.4]
  wire [7:0] _T_25782; // @[Mux.scala 19:72:@20239.4]
  wire [15:0] _T_25783; // @[Mux.scala 19:72:@20240.4]
  wire [15:0] _T_25785; // @[Mux.scala 19:72:@20241.4]
  wire [7:0] _T_25792; // @[Mux.scala 19:72:@20248.4]
  wire [7:0] _T_25799; // @[Mux.scala 19:72:@20255.4]
  wire [15:0] _T_25800; // @[Mux.scala 19:72:@20256.4]
  wire [15:0] _T_25802; // @[Mux.scala 19:72:@20257.4]
  wire [7:0] _T_25809; // @[Mux.scala 19:72:@20264.4]
  wire [7:0] _T_25816; // @[Mux.scala 19:72:@20271.4]
  wire [15:0] _T_25817; // @[Mux.scala 19:72:@20272.4]
  wire [15:0] _T_25819; // @[Mux.scala 19:72:@20273.4]
  wire [7:0] _T_25826; // @[Mux.scala 19:72:@20280.4]
  wire [7:0] _T_25833; // @[Mux.scala 19:72:@20287.4]
  wire [15:0] _T_25834; // @[Mux.scala 19:72:@20288.4]
  wire [15:0] _T_25836; // @[Mux.scala 19:72:@20289.4]
  wire [7:0] _T_25843; // @[Mux.scala 19:72:@20296.4]
  wire [7:0] _T_25850; // @[Mux.scala 19:72:@20303.4]
  wire [15:0] _T_25851; // @[Mux.scala 19:72:@20304.4]
  wire [15:0] _T_25853; // @[Mux.scala 19:72:@20305.4]
  wire [15:0] _T_25868; // @[Mux.scala 19:72:@20320.4]
  wire [15:0] _T_25870; // @[Mux.scala 19:72:@20321.4]
  wire [15:0] _T_25885; // @[Mux.scala 19:72:@20336.4]
  wire [15:0] _T_25887; // @[Mux.scala 19:72:@20337.4]
  wire [15:0] _T_25902; // @[Mux.scala 19:72:@20352.4]
  wire [15:0] _T_25904; // @[Mux.scala 19:72:@20353.4]
  wire [15:0] _T_25919; // @[Mux.scala 19:72:@20368.4]
  wire [15:0] _T_25921; // @[Mux.scala 19:72:@20369.4]
  wire [15:0] _T_25936; // @[Mux.scala 19:72:@20384.4]
  wire [15:0] _T_25938; // @[Mux.scala 19:72:@20385.4]
  wire [15:0] _T_25953; // @[Mux.scala 19:72:@20400.4]
  wire [15:0] _T_25955; // @[Mux.scala 19:72:@20401.4]
  wire [15:0] _T_25970; // @[Mux.scala 19:72:@20416.4]
  wire [15:0] _T_25972; // @[Mux.scala 19:72:@20417.4]
  wire [15:0] _T_25987; // @[Mux.scala 19:72:@20432.4]
  wire [15:0] _T_25989; // @[Mux.scala 19:72:@20433.4]
  wire [15:0] _T_25990; // @[Mux.scala 19:72:@20434.4]
  wire [15:0] _T_25991; // @[Mux.scala 19:72:@20435.4]
  wire [15:0] _T_25992; // @[Mux.scala 19:72:@20436.4]
  wire [15:0] _T_25993; // @[Mux.scala 19:72:@20437.4]
  wire [15:0] _T_25994; // @[Mux.scala 19:72:@20438.4]
  wire [15:0] _T_25995; // @[Mux.scala 19:72:@20439.4]
  wire [15:0] _T_25996; // @[Mux.scala 19:72:@20440.4]
  wire [15:0] _T_25997; // @[Mux.scala 19:72:@20441.4]
  wire [15:0] _T_25998; // @[Mux.scala 19:72:@20442.4]
  wire [15:0] _T_25999; // @[Mux.scala 19:72:@20443.4]
  wire [15:0] _T_26000; // @[Mux.scala 19:72:@20444.4]
  wire [15:0] _T_26001; // @[Mux.scala 19:72:@20445.4]
  wire [15:0] _T_26002; // @[Mux.scala 19:72:@20446.4]
  wire [15:0] _T_26003; // @[Mux.scala 19:72:@20447.4]
  wire [15:0] _T_26004; // @[Mux.scala 19:72:@20448.4]
  wire [7:0] _T_26582; // @[Mux.scala 19:72:@20798.4]
  wire [7:0] _T_26589; // @[Mux.scala 19:72:@20805.4]
  wire [15:0] _T_26590; // @[Mux.scala 19:72:@20806.4]
  wire [15:0] _T_26592; // @[Mux.scala 19:72:@20807.4]
  wire [7:0] _T_26599; // @[Mux.scala 19:72:@20814.4]
  wire [7:0] _T_26606; // @[Mux.scala 19:72:@20821.4]
  wire [15:0] _T_26607; // @[Mux.scala 19:72:@20822.4]
  wire [15:0] _T_26609; // @[Mux.scala 19:72:@20823.4]
  wire [7:0] _T_26616; // @[Mux.scala 19:72:@20830.4]
  wire [7:0] _T_26623; // @[Mux.scala 19:72:@20837.4]
  wire [15:0] _T_26624; // @[Mux.scala 19:72:@20838.4]
  wire [15:0] _T_26626; // @[Mux.scala 19:72:@20839.4]
  wire [7:0] _T_26633; // @[Mux.scala 19:72:@20846.4]
  wire [7:0] _T_26640; // @[Mux.scala 19:72:@20853.4]
  wire [15:0] _T_26641; // @[Mux.scala 19:72:@20854.4]
  wire [15:0] _T_26643; // @[Mux.scala 19:72:@20855.4]
  wire [7:0] _T_26650; // @[Mux.scala 19:72:@20862.4]
  wire [7:0] _T_26657; // @[Mux.scala 19:72:@20869.4]
  wire [15:0] _T_26658; // @[Mux.scala 19:72:@20870.4]
  wire [15:0] _T_26660; // @[Mux.scala 19:72:@20871.4]
  wire [7:0] _T_26667; // @[Mux.scala 19:72:@20878.4]
  wire [7:0] _T_26674; // @[Mux.scala 19:72:@20885.4]
  wire [15:0] _T_26675; // @[Mux.scala 19:72:@20886.4]
  wire [15:0] _T_26677; // @[Mux.scala 19:72:@20887.4]
  wire [7:0] _T_26684; // @[Mux.scala 19:72:@20894.4]
  wire [7:0] _T_26691; // @[Mux.scala 19:72:@20901.4]
  wire [15:0] _T_26692; // @[Mux.scala 19:72:@20902.4]
  wire [15:0] _T_26694; // @[Mux.scala 19:72:@20903.4]
  wire [7:0] _T_26701; // @[Mux.scala 19:72:@20910.4]
  wire [7:0] _T_26708; // @[Mux.scala 19:72:@20917.4]
  wire [15:0] _T_26709; // @[Mux.scala 19:72:@20918.4]
  wire [15:0] _T_26711; // @[Mux.scala 19:72:@20919.4]
  wire [15:0] _T_26726; // @[Mux.scala 19:72:@20934.4]
  wire [15:0] _T_26728; // @[Mux.scala 19:72:@20935.4]
  wire [15:0] _T_26743; // @[Mux.scala 19:72:@20950.4]
  wire [15:0] _T_26745; // @[Mux.scala 19:72:@20951.4]
  wire [15:0] _T_26760; // @[Mux.scala 19:72:@20966.4]
  wire [15:0] _T_26762; // @[Mux.scala 19:72:@20967.4]
  wire [15:0] _T_26777; // @[Mux.scala 19:72:@20982.4]
  wire [15:0] _T_26779; // @[Mux.scala 19:72:@20983.4]
  wire [15:0] _T_26794; // @[Mux.scala 19:72:@20998.4]
  wire [15:0] _T_26796; // @[Mux.scala 19:72:@20999.4]
  wire [15:0] _T_26811; // @[Mux.scala 19:72:@21014.4]
  wire [15:0] _T_26813; // @[Mux.scala 19:72:@21015.4]
  wire [15:0] _T_26828; // @[Mux.scala 19:72:@21030.4]
  wire [15:0] _T_26830; // @[Mux.scala 19:72:@21031.4]
  wire [15:0] _T_26845; // @[Mux.scala 19:72:@21046.4]
  wire [15:0] _T_26847; // @[Mux.scala 19:72:@21047.4]
  wire [15:0] _T_26848; // @[Mux.scala 19:72:@21048.4]
  wire [15:0] _T_26849; // @[Mux.scala 19:72:@21049.4]
  wire [15:0] _T_26850; // @[Mux.scala 19:72:@21050.4]
  wire [15:0] _T_26851; // @[Mux.scala 19:72:@21051.4]
  wire [15:0] _T_26852; // @[Mux.scala 19:72:@21052.4]
  wire [15:0] _T_26853; // @[Mux.scala 19:72:@21053.4]
  wire [15:0] _T_26854; // @[Mux.scala 19:72:@21054.4]
  wire [15:0] _T_26855; // @[Mux.scala 19:72:@21055.4]
  wire [15:0] _T_26856; // @[Mux.scala 19:72:@21056.4]
  wire [15:0] _T_26857; // @[Mux.scala 19:72:@21057.4]
  wire [15:0] _T_26858; // @[Mux.scala 19:72:@21058.4]
  wire [15:0] _T_26859; // @[Mux.scala 19:72:@21059.4]
  wire [15:0] _T_26860; // @[Mux.scala 19:72:@21060.4]
  wire [15:0] _T_26861; // @[Mux.scala 19:72:@21061.4]
  wire [15:0] _T_26862; // @[Mux.scala 19:72:@21062.4]
  wire [7:0] _T_27440; // @[Mux.scala 19:72:@21412.4]
  wire [7:0] _T_27447; // @[Mux.scala 19:72:@21419.4]
  wire [15:0] _T_27448; // @[Mux.scala 19:72:@21420.4]
  wire [15:0] _T_27450; // @[Mux.scala 19:72:@21421.4]
  wire [7:0] _T_27457; // @[Mux.scala 19:72:@21428.4]
  wire [7:0] _T_27464; // @[Mux.scala 19:72:@21435.4]
  wire [15:0] _T_27465; // @[Mux.scala 19:72:@21436.4]
  wire [15:0] _T_27467; // @[Mux.scala 19:72:@21437.4]
  wire [7:0] _T_27474; // @[Mux.scala 19:72:@21444.4]
  wire [7:0] _T_27481; // @[Mux.scala 19:72:@21451.4]
  wire [15:0] _T_27482; // @[Mux.scala 19:72:@21452.4]
  wire [15:0] _T_27484; // @[Mux.scala 19:72:@21453.4]
  wire [7:0] _T_27491; // @[Mux.scala 19:72:@21460.4]
  wire [7:0] _T_27498; // @[Mux.scala 19:72:@21467.4]
  wire [15:0] _T_27499; // @[Mux.scala 19:72:@21468.4]
  wire [15:0] _T_27501; // @[Mux.scala 19:72:@21469.4]
  wire [7:0] _T_27508; // @[Mux.scala 19:72:@21476.4]
  wire [7:0] _T_27515; // @[Mux.scala 19:72:@21483.4]
  wire [15:0] _T_27516; // @[Mux.scala 19:72:@21484.4]
  wire [15:0] _T_27518; // @[Mux.scala 19:72:@21485.4]
  wire [7:0] _T_27525; // @[Mux.scala 19:72:@21492.4]
  wire [7:0] _T_27532; // @[Mux.scala 19:72:@21499.4]
  wire [15:0] _T_27533; // @[Mux.scala 19:72:@21500.4]
  wire [15:0] _T_27535; // @[Mux.scala 19:72:@21501.4]
  wire [7:0] _T_27542; // @[Mux.scala 19:72:@21508.4]
  wire [7:0] _T_27549; // @[Mux.scala 19:72:@21515.4]
  wire [15:0] _T_27550; // @[Mux.scala 19:72:@21516.4]
  wire [15:0] _T_27552; // @[Mux.scala 19:72:@21517.4]
  wire [7:0] _T_27559; // @[Mux.scala 19:72:@21524.4]
  wire [7:0] _T_27566; // @[Mux.scala 19:72:@21531.4]
  wire [15:0] _T_27567; // @[Mux.scala 19:72:@21532.4]
  wire [15:0] _T_27569; // @[Mux.scala 19:72:@21533.4]
  wire [15:0] _T_27584; // @[Mux.scala 19:72:@21548.4]
  wire [15:0] _T_27586; // @[Mux.scala 19:72:@21549.4]
  wire [15:0] _T_27601; // @[Mux.scala 19:72:@21564.4]
  wire [15:0] _T_27603; // @[Mux.scala 19:72:@21565.4]
  wire [15:0] _T_27618; // @[Mux.scala 19:72:@21580.4]
  wire [15:0] _T_27620; // @[Mux.scala 19:72:@21581.4]
  wire [15:0] _T_27635; // @[Mux.scala 19:72:@21596.4]
  wire [15:0] _T_27637; // @[Mux.scala 19:72:@21597.4]
  wire [15:0] _T_27652; // @[Mux.scala 19:72:@21612.4]
  wire [15:0] _T_27654; // @[Mux.scala 19:72:@21613.4]
  wire [15:0] _T_27669; // @[Mux.scala 19:72:@21628.4]
  wire [15:0] _T_27671; // @[Mux.scala 19:72:@21629.4]
  wire [15:0] _T_27686; // @[Mux.scala 19:72:@21644.4]
  wire [15:0] _T_27688; // @[Mux.scala 19:72:@21645.4]
  wire [15:0] _T_27703; // @[Mux.scala 19:72:@21660.4]
  wire [15:0] _T_27705; // @[Mux.scala 19:72:@21661.4]
  wire [15:0] _T_27706; // @[Mux.scala 19:72:@21662.4]
  wire [15:0] _T_27707; // @[Mux.scala 19:72:@21663.4]
  wire [15:0] _T_27708; // @[Mux.scala 19:72:@21664.4]
  wire [15:0] _T_27709; // @[Mux.scala 19:72:@21665.4]
  wire [15:0] _T_27710; // @[Mux.scala 19:72:@21666.4]
  wire [15:0] _T_27711; // @[Mux.scala 19:72:@21667.4]
  wire [15:0] _T_27712; // @[Mux.scala 19:72:@21668.4]
  wire [15:0] _T_27713; // @[Mux.scala 19:72:@21669.4]
  wire [15:0] _T_27714; // @[Mux.scala 19:72:@21670.4]
  wire [15:0] _T_27715; // @[Mux.scala 19:72:@21671.4]
  wire [15:0] _T_27716; // @[Mux.scala 19:72:@21672.4]
  wire [15:0] _T_27717; // @[Mux.scala 19:72:@21673.4]
  wire [15:0] _T_27718; // @[Mux.scala 19:72:@21674.4]
  wire [15:0] _T_27719; // @[Mux.scala 19:72:@21675.4]
  wire [15:0] _T_27720; // @[Mux.scala 19:72:@21676.4]
  wire [7:0] _T_28298; // @[Mux.scala 19:72:@22026.4]
  wire [7:0] _T_28305; // @[Mux.scala 19:72:@22033.4]
  wire [15:0] _T_28306; // @[Mux.scala 19:72:@22034.4]
  wire [15:0] _T_28308; // @[Mux.scala 19:72:@22035.4]
  wire [7:0] _T_28315; // @[Mux.scala 19:72:@22042.4]
  wire [7:0] _T_28322; // @[Mux.scala 19:72:@22049.4]
  wire [15:0] _T_28323; // @[Mux.scala 19:72:@22050.4]
  wire [15:0] _T_28325; // @[Mux.scala 19:72:@22051.4]
  wire [7:0] _T_28332; // @[Mux.scala 19:72:@22058.4]
  wire [7:0] _T_28339; // @[Mux.scala 19:72:@22065.4]
  wire [15:0] _T_28340; // @[Mux.scala 19:72:@22066.4]
  wire [15:0] _T_28342; // @[Mux.scala 19:72:@22067.4]
  wire [7:0] _T_28349; // @[Mux.scala 19:72:@22074.4]
  wire [7:0] _T_28356; // @[Mux.scala 19:72:@22081.4]
  wire [15:0] _T_28357; // @[Mux.scala 19:72:@22082.4]
  wire [15:0] _T_28359; // @[Mux.scala 19:72:@22083.4]
  wire [7:0] _T_28366; // @[Mux.scala 19:72:@22090.4]
  wire [7:0] _T_28373; // @[Mux.scala 19:72:@22097.4]
  wire [15:0] _T_28374; // @[Mux.scala 19:72:@22098.4]
  wire [15:0] _T_28376; // @[Mux.scala 19:72:@22099.4]
  wire [7:0] _T_28383; // @[Mux.scala 19:72:@22106.4]
  wire [7:0] _T_28390; // @[Mux.scala 19:72:@22113.4]
  wire [15:0] _T_28391; // @[Mux.scala 19:72:@22114.4]
  wire [15:0] _T_28393; // @[Mux.scala 19:72:@22115.4]
  wire [7:0] _T_28400; // @[Mux.scala 19:72:@22122.4]
  wire [7:0] _T_28407; // @[Mux.scala 19:72:@22129.4]
  wire [15:0] _T_28408; // @[Mux.scala 19:72:@22130.4]
  wire [15:0] _T_28410; // @[Mux.scala 19:72:@22131.4]
  wire [7:0] _T_28417; // @[Mux.scala 19:72:@22138.4]
  wire [7:0] _T_28424; // @[Mux.scala 19:72:@22145.4]
  wire [15:0] _T_28425; // @[Mux.scala 19:72:@22146.4]
  wire [15:0] _T_28427; // @[Mux.scala 19:72:@22147.4]
  wire [15:0] _T_28442; // @[Mux.scala 19:72:@22162.4]
  wire [15:0] _T_28444; // @[Mux.scala 19:72:@22163.4]
  wire [15:0] _T_28459; // @[Mux.scala 19:72:@22178.4]
  wire [15:0] _T_28461; // @[Mux.scala 19:72:@22179.4]
  wire [15:0] _T_28476; // @[Mux.scala 19:72:@22194.4]
  wire [15:0] _T_28478; // @[Mux.scala 19:72:@22195.4]
  wire [15:0] _T_28493; // @[Mux.scala 19:72:@22210.4]
  wire [15:0] _T_28495; // @[Mux.scala 19:72:@22211.4]
  wire [15:0] _T_28510; // @[Mux.scala 19:72:@22226.4]
  wire [15:0] _T_28512; // @[Mux.scala 19:72:@22227.4]
  wire [15:0] _T_28527; // @[Mux.scala 19:72:@22242.4]
  wire [15:0] _T_28529; // @[Mux.scala 19:72:@22243.4]
  wire [15:0] _T_28544; // @[Mux.scala 19:72:@22258.4]
  wire [15:0] _T_28546; // @[Mux.scala 19:72:@22259.4]
  wire [15:0] _T_28561; // @[Mux.scala 19:72:@22274.4]
  wire [15:0] _T_28563; // @[Mux.scala 19:72:@22275.4]
  wire [15:0] _T_28564; // @[Mux.scala 19:72:@22276.4]
  wire [15:0] _T_28565; // @[Mux.scala 19:72:@22277.4]
  wire [15:0] _T_28566; // @[Mux.scala 19:72:@22278.4]
  wire [15:0] _T_28567; // @[Mux.scala 19:72:@22279.4]
  wire [15:0] _T_28568; // @[Mux.scala 19:72:@22280.4]
  wire [15:0] _T_28569; // @[Mux.scala 19:72:@22281.4]
  wire [15:0] _T_28570; // @[Mux.scala 19:72:@22282.4]
  wire [15:0] _T_28571; // @[Mux.scala 19:72:@22283.4]
  wire [15:0] _T_28572; // @[Mux.scala 19:72:@22284.4]
  wire [15:0] _T_28573; // @[Mux.scala 19:72:@22285.4]
  wire [15:0] _T_28574; // @[Mux.scala 19:72:@22286.4]
  wire [15:0] _T_28575; // @[Mux.scala 19:72:@22287.4]
  wire [15:0] _T_28576; // @[Mux.scala 19:72:@22288.4]
  wire [15:0] _T_28577; // @[Mux.scala 19:72:@22289.4]
  wire [15:0] _T_28578; // @[Mux.scala 19:72:@22290.4]
  wire [7:0] _T_29156; // @[Mux.scala 19:72:@22640.4]
  wire [7:0] _T_29163; // @[Mux.scala 19:72:@22647.4]
  wire [15:0] _T_29164; // @[Mux.scala 19:72:@22648.4]
  wire [15:0] _T_29166; // @[Mux.scala 19:72:@22649.4]
  wire [7:0] _T_29173; // @[Mux.scala 19:72:@22656.4]
  wire [7:0] _T_29180; // @[Mux.scala 19:72:@22663.4]
  wire [15:0] _T_29181; // @[Mux.scala 19:72:@22664.4]
  wire [15:0] _T_29183; // @[Mux.scala 19:72:@22665.4]
  wire [7:0] _T_29190; // @[Mux.scala 19:72:@22672.4]
  wire [7:0] _T_29197; // @[Mux.scala 19:72:@22679.4]
  wire [15:0] _T_29198; // @[Mux.scala 19:72:@22680.4]
  wire [15:0] _T_29200; // @[Mux.scala 19:72:@22681.4]
  wire [7:0] _T_29207; // @[Mux.scala 19:72:@22688.4]
  wire [7:0] _T_29214; // @[Mux.scala 19:72:@22695.4]
  wire [15:0] _T_29215; // @[Mux.scala 19:72:@22696.4]
  wire [15:0] _T_29217; // @[Mux.scala 19:72:@22697.4]
  wire [7:0] _T_29224; // @[Mux.scala 19:72:@22704.4]
  wire [7:0] _T_29231; // @[Mux.scala 19:72:@22711.4]
  wire [15:0] _T_29232; // @[Mux.scala 19:72:@22712.4]
  wire [15:0] _T_29234; // @[Mux.scala 19:72:@22713.4]
  wire [7:0] _T_29241; // @[Mux.scala 19:72:@22720.4]
  wire [7:0] _T_29248; // @[Mux.scala 19:72:@22727.4]
  wire [15:0] _T_29249; // @[Mux.scala 19:72:@22728.4]
  wire [15:0] _T_29251; // @[Mux.scala 19:72:@22729.4]
  wire [7:0] _T_29258; // @[Mux.scala 19:72:@22736.4]
  wire [7:0] _T_29265; // @[Mux.scala 19:72:@22743.4]
  wire [15:0] _T_29266; // @[Mux.scala 19:72:@22744.4]
  wire [15:0] _T_29268; // @[Mux.scala 19:72:@22745.4]
  wire [7:0] _T_29275; // @[Mux.scala 19:72:@22752.4]
  wire [7:0] _T_29282; // @[Mux.scala 19:72:@22759.4]
  wire [15:0] _T_29283; // @[Mux.scala 19:72:@22760.4]
  wire [15:0] _T_29285; // @[Mux.scala 19:72:@22761.4]
  wire [15:0] _T_29300; // @[Mux.scala 19:72:@22776.4]
  wire [15:0] _T_29302; // @[Mux.scala 19:72:@22777.4]
  wire [15:0] _T_29317; // @[Mux.scala 19:72:@22792.4]
  wire [15:0] _T_29319; // @[Mux.scala 19:72:@22793.4]
  wire [15:0] _T_29334; // @[Mux.scala 19:72:@22808.4]
  wire [15:0] _T_29336; // @[Mux.scala 19:72:@22809.4]
  wire [15:0] _T_29351; // @[Mux.scala 19:72:@22824.4]
  wire [15:0] _T_29353; // @[Mux.scala 19:72:@22825.4]
  wire [15:0] _T_29368; // @[Mux.scala 19:72:@22840.4]
  wire [15:0] _T_29370; // @[Mux.scala 19:72:@22841.4]
  wire [15:0] _T_29385; // @[Mux.scala 19:72:@22856.4]
  wire [15:0] _T_29387; // @[Mux.scala 19:72:@22857.4]
  wire [15:0] _T_29402; // @[Mux.scala 19:72:@22872.4]
  wire [15:0] _T_29404; // @[Mux.scala 19:72:@22873.4]
  wire [15:0] _T_29419; // @[Mux.scala 19:72:@22888.4]
  wire [15:0] _T_29421; // @[Mux.scala 19:72:@22889.4]
  wire [15:0] _T_29422; // @[Mux.scala 19:72:@22890.4]
  wire [15:0] _T_29423; // @[Mux.scala 19:72:@22891.4]
  wire [15:0] _T_29424; // @[Mux.scala 19:72:@22892.4]
  wire [15:0] _T_29425; // @[Mux.scala 19:72:@22893.4]
  wire [15:0] _T_29426; // @[Mux.scala 19:72:@22894.4]
  wire [15:0] _T_29427; // @[Mux.scala 19:72:@22895.4]
  wire [15:0] _T_29428; // @[Mux.scala 19:72:@22896.4]
  wire [15:0] _T_29429; // @[Mux.scala 19:72:@22897.4]
  wire [15:0] _T_29430; // @[Mux.scala 19:72:@22898.4]
  wire [15:0] _T_29431; // @[Mux.scala 19:72:@22899.4]
  wire [15:0] _T_29432; // @[Mux.scala 19:72:@22900.4]
  wire [15:0] _T_29433; // @[Mux.scala 19:72:@22901.4]
  wire [15:0] _T_29434; // @[Mux.scala 19:72:@22902.4]
  wire [15:0] _T_29435; // @[Mux.scala 19:72:@22903.4]
  wire [15:0] _T_29436; // @[Mux.scala 19:72:@22904.4]
  wire [7:0] _T_30014; // @[Mux.scala 19:72:@23254.4]
  wire [7:0] _T_30021; // @[Mux.scala 19:72:@23261.4]
  wire [15:0] _T_30022; // @[Mux.scala 19:72:@23262.4]
  wire [15:0] _T_30024; // @[Mux.scala 19:72:@23263.4]
  wire [7:0] _T_30031; // @[Mux.scala 19:72:@23270.4]
  wire [7:0] _T_30038; // @[Mux.scala 19:72:@23277.4]
  wire [15:0] _T_30039; // @[Mux.scala 19:72:@23278.4]
  wire [15:0] _T_30041; // @[Mux.scala 19:72:@23279.4]
  wire [7:0] _T_30048; // @[Mux.scala 19:72:@23286.4]
  wire [7:0] _T_30055; // @[Mux.scala 19:72:@23293.4]
  wire [15:0] _T_30056; // @[Mux.scala 19:72:@23294.4]
  wire [15:0] _T_30058; // @[Mux.scala 19:72:@23295.4]
  wire [7:0] _T_30065; // @[Mux.scala 19:72:@23302.4]
  wire [7:0] _T_30072; // @[Mux.scala 19:72:@23309.4]
  wire [15:0] _T_30073; // @[Mux.scala 19:72:@23310.4]
  wire [15:0] _T_30075; // @[Mux.scala 19:72:@23311.4]
  wire [7:0] _T_30082; // @[Mux.scala 19:72:@23318.4]
  wire [7:0] _T_30089; // @[Mux.scala 19:72:@23325.4]
  wire [15:0] _T_30090; // @[Mux.scala 19:72:@23326.4]
  wire [15:0] _T_30092; // @[Mux.scala 19:72:@23327.4]
  wire [7:0] _T_30099; // @[Mux.scala 19:72:@23334.4]
  wire [7:0] _T_30106; // @[Mux.scala 19:72:@23341.4]
  wire [15:0] _T_30107; // @[Mux.scala 19:72:@23342.4]
  wire [15:0] _T_30109; // @[Mux.scala 19:72:@23343.4]
  wire [7:0] _T_30116; // @[Mux.scala 19:72:@23350.4]
  wire [7:0] _T_30123; // @[Mux.scala 19:72:@23357.4]
  wire [15:0] _T_30124; // @[Mux.scala 19:72:@23358.4]
  wire [15:0] _T_30126; // @[Mux.scala 19:72:@23359.4]
  wire [7:0] _T_30133; // @[Mux.scala 19:72:@23366.4]
  wire [7:0] _T_30140; // @[Mux.scala 19:72:@23373.4]
  wire [15:0] _T_30141; // @[Mux.scala 19:72:@23374.4]
  wire [15:0] _T_30143; // @[Mux.scala 19:72:@23375.4]
  wire [15:0] _T_30158; // @[Mux.scala 19:72:@23390.4]
  wire [15:0] _T_30160; // @[Mux.scala 19:72:@23391.4]
  wire [15:0] _T_30175; // @[Mux.scala 19:72:@23406.4]
  wire [15:0] _T_30177; // @[Mux.scala 19:72:@23407.4]
  wire [15:0] _T_30192; // @[Mux.scala 19:72:@23422.4]
  wire [15:0] _T_30194; // @[Mux.scala 19:72:@23423.4]
  wire [15:0] _T_30209; // @[Mux.scala 19:72:@23438.4]
  wire [15:0] _T_30211; // @[Mux.scala 19:72:@23439.4]
  wire [15:0] _T_30226; // @[Mux.scala 19:72:@23454.4]
  wire [15:0] _T_30228; // @[Mux.scala 19:72:@23455.4]
  wire [15:0] _T_30243; // @[Mux.scala 19:72:@23470.4]
  wire [15:0] _T_30245; // @[Mux.scala 19:72:@23471.4]
  wire [15:0] _T_30260; // @[Mux.scala 19:72:@23486.4]
  wire [15:0] _T_30262; // @[Mux.scala 19:72:@23487.4]
  wire [15:0] _T_30277; // @[Mux.scala 19:72:@23502.4]
  wire [15:0] _T_30279; // @[Mux.scala 19:72:@23503.4]
  wire [15:0] _T_30280; // @[Mux.scala 19:72:@23504.4]
  wire [15:0] _T_30281; // @[Mux.scala 19:72:@23505.4]
  wire [15:0] _T_30282; // @[Mux.scala 19:72:@23506.4]
  wire [15:0] _T_30283; // @[Mux.scala 19:72:@23507.4]
  wire [15:0] _T_30284; // @[Mux.scala 19:72:@23508.4]
  wire [15:0] _T_30285; // @[Mux.scala 19:72:@23509.4]
  wire [15:0] _T_30286; // @[Mux.scala 19:72:@23510.4]
  wire [15:0] _T_30287; // @[Mux.scala 19:72:@23511.4]
  wire [15:0] _T_30288; // @[Mux.scala 19:72:@23512.4]
  wire [15:0] _T_30289; // @[Mux.scala 19:72:@23513.4]
  wire [15:0] _T_30290; // @[Mux.scala 19:72:@23514.4]
  wire [15:0] _T_30291; // @[Mux.scala 19:72:@23515.4]
  wire [15:0] _T_30292; // @[Mux.scala 19:72:@23516.4]
  wire [15:0] _T_30293; // @[Mux.scala 19:72:@23517.4]
  wire [15:0] _T_30294; // @[Mux.scala 19:72:@23518.4]
  wire [7:0] _T_30872; // @[Mux.scala 19:72:@23868.4]
  wire [7:0] _T_30879; // @[Mux.scala 19:72:@23875.4]
  wire [15:0] _T_30880; // @[Mux.scala 19:72:@23876.4]
  wire [15:0] _T_30882; // @[Mux.scala 19:72:@23877.4]
  wire [7:0] _T_30889; // @[Mux.scala 19:72:@23884.4]
  wire [7:0] _T_30896; // @[Mux.scala 19:72:@23891.4]
  wire [15:0] _T_30897; // @[Mux.scala 19:72:@23892.4]
  wire [15:0] _T_30899; // @[Mux.scala 19:72:@23893.4]
  wire [7:0] _T_30906; // @[Mux.scala 19:72:@23900.4]
  wire [7:0] _T_30913; // @[Mux.scala 19:72:@23907.4]
  wire [15:0] _T_30914; // @[Mux.scala 19:72:@23908.4]
  wire [15:0] _T_30916; // @[Mux.scala 19:72:@23909.4]
  wire [7:0] _T_30923; // @[Mux.scala 19:72:@23916.4]
  wire [7:0] _T_30930; // @[Mux.scala 19:72:@23923.4]
  wire [15:0] _T_30931; // @[Mux.scala 19:72:@23924.4]
  wire [15:0] _T_30933; // @[Mux.scala 19:72:@23925.4]
  wire [7:0] _T_30940; // @[Mux.scala 19:72:@23932.4]
  wire [7:0] _T_30947; // @[Mux.scala 19:72:@23939.4]
  wire [15:0] _T_30948; // @[Mux.scala 19:72:@23940.4]
  wire [15:0] _T_30950; // @[Mux.scala 19:72:@23941.4]
  wire [7:0] _T_30957; // @[Mux.scala 19:72:@23948.4]
  wire [7:0] _T_30964; // @[Mux.scala 19:72:@23955.4]
  wire [15:0] _T_30965; // @[Mux.scala 19:72:@23956.4]
  wire [15:0] _T_30967; // @[Mux.scala 19:72:@23957.4]
  wire [7:0] _T_30974; // @[Mux.scala 19:72:@23964.4]
  wire [7:0] _T_30981; // @[Mux.scala 19:72:@23971.4]
  wire [15:0] _T_30982; // @[Mux.scala 19:72:@23972.4]
  wire [15:0] _T_30984; // @[Mux.scala 19:72:@23973.4]
  wire [7:0] _T_30991; // @[Mux.scala 19:72:@23980.4]
  wire [7:0] _T_30998; // @[Mux.scala 19:72:@23987.4]
  wire [15:0] _T_30999; // @[Mux.scala 19:72:@23988.4]
  wire [15:0] _T_31001; // @[Mux.scala 19:72:@23989.4]
  wire [15:0] _T_31016; // @[Mux.scala 19:72:@24004.4]
  wire [15:0] _T_31018; // @[Mux.scala 19:72:@24005.4]
  wire [15:0] _T_31033; // @[Mux.scala 19:72:@24020.4]
  wire [15:0] _T_31035; // @[Mux.scala 19:72:@24021.4]
  wire [15:0] _T_31050; // @[Mux.scala 19:72:@24036.4]
  wire [15:0] _T_31052; // @[Mux.scala 19:72:@24037.4]
  wire [15:0] _T_31067; // @[Mux.scala 19:72:@24052.4]
  wire [15:0] _T_31069; // @[Mux.scala 19:72:@24053.4]
  wire [15:0] _T_31084; // @[Mux.scala 19:72:@24068.4]
  wire [15:0] _T_31086; // @[Mux.scala 19:72:@24069.4]
  wire [15:0] _T_31101; // @[Mux.scala 19:72:@24084.4]
  wire [15:0] _T_31103; // @[Mux.scala 19:72:@24085.4]
  wire [15:0] _T_31118; // @[Mux.scala 19:72:@24100.4]
  wire [15:0] _T_31120; // @[Mux.scala 19:72:@24101.4]
  wire [15:0] _T_31135; // @[Mux.scala 19:72:@24116.4]
  wire [15:0] _T_31137; // @[Mux.scala 19:72:@24117.4]
  wire [15:0] _T_31138; // @[Mux.scala 19:72:@24118.4]
  wire [15:0] _T_31139; // @[Mux.scala 19:72:@24119.4]
  wire [15:0] _T_31140; // @[Mux.scala 19:72:@24120.4]
  wire [15:0] _T_31141; // @[Mux.scala 19:72:@24121.4]
  wire [15:0] _T_31142; // @[Mux.scala 19:72:@24122.4]
  wire [15:0] _T_31143; // @[Mux.scala 19:72:@24123.4]
  wire [15:0] _T_31144; // @[Mux.scala 19:72:@24124.4]
  wire [15:0] _T_31145; // @[Mux.scala 19:72:@24125.4]
  wire [15:0] _T_31146; // @[Mux.scala 19:72:@24126.4]
  wire [15:0] _T_31147; // @[Mux.scala 19:72:@24127.4]
  wire [15:0] _T_31148; // @[Mux.scala 19:72:@24128.4]
  wire [15:0] _T_31149; // @[Mux.scala 19:72:@24129.4]
  wire [15:0] _T_31150; // @[Mux.scala 19:72:@24130.4]
  wire [15:0] _T_31151; // @[Mux.scala 19:72:@24131.4]
  wire [15:0] _T_31152; // @[Mux.scala 19:72:@24132.4]
  reg  conflictPReg_0_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_163;
  reg  conflictPReg_0_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_164;
  reg  conflictPReg_0_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_165;
  reg  conflictPReg_0_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_166;
  reg  conflictPReg_0_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_167;
  reg  conflictPReg_0_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_168;
  reg  conflictPReg_0_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_169;
  reg  conflictPReg_0_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_170;
  reg  conflictPReg_0_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_171;
  reg  conflictPReg_0_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_172;
  reg  conflictPReg_0_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_173;
  reg  conflictPReg_0_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_174;
  reg  conflictPReg_0_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_175;
  reg  conflictPReg_0_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_176;
  reg  conflictPReg_0_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_177;
  reg  conflictPReg_0_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_178;
  reg  conflictPReg_1_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_179;
  reg  conflictPReg_1_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_180;
  reg  conflictPReg_1_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_181;
  reg  conflictPReg_1_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_182;
  reg  conflictPReg_1_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_183;
  reg  conflictPReg_1_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_184;
  reg  conflictPReg_1_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_185;
  reg  conflictPReg_1_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_186;
  reg  conflictPReg_1_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_187;
  reg  conflictPReg_1_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_188;
  reg  conflictPReg_1_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_189;
  reg  conflictPReg_1_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_190;
  reg  conflictPReg_1_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_191;
  reg  conflictPReg_1_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_192;
  reg  conflictPReg_1_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_193;
  reg  conflictPReg_1_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_194;
  reg  conflictPReg_2_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_195;
  reg  conflictPReg_2_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_196;
  reg  conflictPReg_2_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_197;
  reg  conflictPReg_2_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_198;
  reg  conflictPReg_2_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_199;
  reg  conflictPReg_2_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_200;
  reg  conflictPReg_2_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_201;
  reg  conflictPReg_2_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_202;
  reg  conflictPReg_2_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_203;
  reg  conflictPReg_2_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_204;
  reg  conflictPReg_2_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_205;
  reg  conflictPReg_2_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_206;
  reg  conflictPReg_2_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_207;
  reg  conflictPReg_2_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_208;
  reg  conflictPReg_2_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_209;
  reg  conflictPReg_2_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_210;
  reg  conflictPReg_3_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_211;
  reg  conflictPReg_3_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_212;
  reg  conflictPReg_3_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_213;
  reg  conflictPReg_3_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_214;
  reg  conflictPReg_3_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_215;
  reg  conflictPReg_3_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_216;
  reg  conflictPReg_3_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_217;
  reg  conflictPReg_3_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_218;
  reg  conflictPReg_3_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_219;
  reg  conflictPReg_3_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_220;
  reg  conflictPReg_3_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_221;
  reg  conflictPReg_3_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_222;
  reg  conflictPReg_3_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_223;
  reg  conflictPReg_3_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_224;
  reg  conflictPReg_3_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_225;
  reg  conflictPReg_3_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_226;
  reg  conflictPReg_4_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_227;
  reg  conflictPReg_4_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_228;
  reg  conflictPReg_4_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_229;
  reg  conflictPReg_4_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_230;
  reg  conflictPReg_4_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_231;
  reg  conflictPReg_4_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_232;
  reg  conflictPReg_4_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_233;
  reg  conflictPReg_4_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_234;
  reg  conflictPReg_4_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_235;
  reg  conflictPReg_4_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_236;
  reg  conflictPReg_4_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_237;
  reg  conflictPReg_4_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_238;
  reg  conflictPReg_4_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_239;
  reg  conflictPReg_4_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_240;
  reg  conflictPReg_4_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_241;
  reg  conflictPReg_4_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_242;
  reg  conflictPReg_5_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_243;
  reg  conflictPReg_5_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_244;
  reg  conflictPReg_5_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_245;
  reg  conflictPReg_5_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_246;
  reg  conflictPReg_5_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_247;
  reg  conflictPReg_5_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_248;
  reg  conflictPReg_5_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_249;
  reg  conflictPReg_5_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_250;
  reg  conflictPReg_5_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_251;
  reg  conflictPReg_5_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_252;
  reg  conflictPReg_5_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_253;
  reg  conflictPReg_5_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_254;
  reg  conflictPReg_5_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_255;
  reg  conflictPReg_5_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_256;
  reg  conflictPReg_5_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_257;
  reg  conflictPReg_5_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_258;
  reg  conflictPReg_6_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_259;
  reg  conflictPReg_6_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_260;
  reg  conflictPReg_6_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_261;
  reg  conflictPReg_6_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_262;
  reg  conflictPReg_6_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_263;
  reg  conflictPReg_6_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_264;
  reg  conflictPReg_6_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_265;
  reg  conflictPReg_6_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_266;
  reg  conflictPReg_6_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_267;
  reg  conflictPReg_6_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_268;
  reg  conflictPReg_6_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_269;
  reg  conflictPReg_6_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_270;
  reg  conflictPReg_6_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_271;
  reg  conflictPReg_6_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_272;
  reg  conflictPReg_6_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_273;
  reg  conflictPReg_6_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_274;
  reg  conflictPReg_7_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_275;
  reg  conflictPReg_7_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_276;
  reg  conflictPReg_7_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_277;
  reg  conflictPReg_7_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_278;
  reg  conflictPReg_7_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_279;
  reg  conflictPReg_7_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_280;
  reg  conflictPReg_7_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_281;
  reg  conflictPReg_7_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_282;
  reg  conflictPReg_7_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_283;
  reg  conflictPReg_7_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_284;
  reg  conflictPReg_7_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_285;
  reg  conflictPReg_7_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_286;
  reg  conflictPReg_7_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_287;
  reg  conflictPReg_7_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_288;
  reg  conflictPReg_7_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_289;
  reg  conflictPReg_7_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_290;
  reg  conflictPReg_8_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_291;
  reg  conflictPReg_8_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_292;
  reg  conflictPReg_8_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_293;
  reg  conflictPReg_8_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_294;
  reg  conflictPReg_8_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_295;
  reg  conflictPReg_8_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_296;
  reg  conflictPReg_8_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_297;
  reg  conflictPReg_8_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_298;
  reg  conflictPReg_8_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_299;
  reg  conflictPReg_8_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_300;
  reg  conflictPReg_8_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_301;
  reg  conflictPReg_8_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_302;
  reg  conflictPReg_8_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_303;
  reg  conflictPReg_8_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_304;
  reg  conflictPReg_8_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_305;
  reg  conflictPReg_8_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_306;
  reg  conflictPReg_9_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_307;
  reg  conflictPReg_9_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_308;
  reg  conflictPReg_9_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_309;
  reg  conflictPReg_9_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_310;
  reg  conflictPReg_9_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_311;
  reg  conflictPReg_9_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_312;
  reg  conflictPReg_9_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_313;
  reg  conflictPReg_9_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_314;
  reg  conflictPReg_9_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_315;
  reg  conflictPReg_9_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_316;
  reg  conflictPReg_9_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_317;
  reg  conflictPReg_9_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_318;
  reg  conflictPReg_9_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_319;
  reg  conflictPReg_9_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_320;
  reg  conflictPReg_9_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_321;
  reg  conflictPReg_9_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_322;
  reg  conflictPReg_10_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_323;
  reg  conflictPReg_10_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_324;
  reg  conflictPReg_10_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_325;
  reg  conflictPReg_10_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_326;
  reg  conflictPReg_10_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_327;
  reg  conflictPReg_10_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_328;
  reg  conflictPReg_10_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_329;
  reg  conflictPReg_10_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_330;
  reg  conflictPReg_10_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_331;
  reg  conflictPReg_10_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_332;
  reg  conflictPReg_10_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_333;
  reg  conflictPReg_10_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_334;
  reg  conflictPReg_10_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_335;
  reg  conflictPReg_10_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_336;
  reg  conflictPReg_10_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_337;
  reg  conflictPReg_10_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_338;
  reg  conflictPReg_11_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_339;
  reg  conflictPReg_11_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_340;
  reg  conflictPReg_11_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_341;
  reg  conflictPReg_11_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_342;
  reg  conflictPReg_11_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_343;
  reg  conflictPReg_11_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_344;
  reg  conflictPReg_11_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_345;
  reg  conflictPReg_11_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_346;
  reg  conflictPReg_11_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_347;
  reg  conflictPReg_11_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_348;
  reg  conflictPReg_11_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_349;
  reg  conflictPReg_11_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_350;
  reg  conflictPReg_11_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_351;
  reg  conflictPReg_11_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_352;
  reg  conflictPReg_11_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_353;
  reg  conflictPReg_11_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_354;
  reg  conflictPReg_12_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_355;
  reg  conflictPReg_12_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_356;
  reg  conflictPReg_12_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_357;
  reg  conflictPReg_12_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_358;
  reg  conflictPReg_12_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_359;
  reg  conflictPReg_12_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_360;
  reg  conflictPReg_12_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_361;
  reg  conflictPReg_12_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_362;
  reg  conflictPReg_12_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_363;
  reg  conflictPReg_12_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_364;
  reg  conflictPReg_12_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_365;
  reg  conflictPReg_12_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_366;
  reg  conflictPReg_12_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_367;
  reg  conflictPReg_12_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_368;
  reg  conflictPReg_12_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_369;
  reg  conflictPReg_12_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_370;
  reg  conflictPReg_13_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_371;
  reg  conflictPReg_13_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_372;
  reg  conflictPReg_13_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_373;
  reg  conflictPReg_13_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_374;
  reg  conflictPReg_13_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_375;
  reg  conflictPReg_13_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_376;
  reg  conflictPReg_13_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_377;
  reg  conflictPReg_13_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_378;
  reg  conflictPReg_13_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_379;
  reg  conflictPReg_13_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_380;
  reg  conflictPReg_13_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_381;
  reg  conflictPReg_13_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_382;
  reg  conflictPReg_13_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_383;
  reg  conflictPReg_13_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_384;
  reg  conflictPReg_13_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_385;
  reg  conflictPReg_13_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_386;
  reg  conflictPReg_14_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_387;
  reg  conflictPReg_14_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_388;
  reg  conflictPReg_14_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_389;
  reg  conflictPReg_14_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_390;
  reg  conflictPReg_14_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_391;
  reg  conflictPReg_14_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_392;
  reg  conflictPReg_14_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_393;
  reg  conflictPReg_14_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_394;
  reg  conflictPReg_14_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_395;
  reg  conflictPReg_14_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_396;
  reg  conflictPReg_14_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_397;
  reg  conflictPReg_14_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_398;
  reg  conflictPReg_14_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_399;
  reg  conflictPReg_14_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_400;
  reg  conflictPReg_14_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_401;
  reg  conflictPReg_14_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_402;
  reg  conflictPReg_15_0; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_403;
  reg  conflictPReg_15_1; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_404;
  reg  conflictPReg_15_2; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_405;
  reg  conflictPReg_15_3; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_406;
  reg  conflictPReg_15_4; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_407;
  reg  conflictPReg_15_5; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_408;
  reg  conflictPReg_15_6; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_409;
  reg  conflictPReg_15_7; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_410;
  reg  conflictPReg_15_8; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_411;
  reg  conflictPReg_15_9; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_412;
  reg  conflictPReg_15_10; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_413;
  reg  conflictPReg_15_11; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_414;
  reg  conflictPReg_15_12; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_415;
  reg  conflictPReg_15_13; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_416;
  reg  conflictPReg_15_14; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_417;
  reg  conflictPReg_15_15; // @[LoadQueue.scala 166:29:@24425.4]
  reg [31:0] _RAND_418;
  wire [7:0] _T_52326; // @[Mux.scala 19:72:@24996.4]
  wire [7:0] _T_52333; // @[Mux.scala 19:72:@25003.4]
  wire [15:0] _T_52334; // @[Mux.scala 19:72:@25004.4]
  wire [15:0] _T_52336; // @[Mux.scala 19:72:@25005.4]
  wire [7:0] _T_52343; // @[Mux.scala 19:72:@25012.4]
  wire [7:0] _T_52350; // @[Mux.scala 19:72:@25019.4]
  wire [15:0] _T_52351; // @[Mux.scala 19:72:@25020.4]
  wire [15:0] _T_52353; // @[Mux.scala 19:72:@25021.4]
  wire [7:0] _T_52360; // @[Mux.scala 19:72:@25028.4]
  wire [7:0] _T_52367; // @[Mux.scala 19:72:@25035.4]
  wire [15:0] _T_52368; // @[Mux.scala 19:72:@25036.4]
  wire [15:0] _T_52370; // @[Mux.scala 19:72:@25037.4]
  wire [7:0] _T_52377; // @[Mux.scala 19:72:@25044.4]
  wire [7:0] _T_52384; // @[Mux.scala 19:72:@25051.4]
  wire [15:0] _T_52385; // @[Mux.scala 19:72:@25052.4]
  wire [15:0] _T_52387; // @[Mux.scala 19:72:@25053.4]
  wire [7:0] _T_52394; // @[Mux.scala 19:72:@25060.4]
  wire [7:0] _T_52401; // @[Mux.scala 19:72:@25067.4]
  wire [15:0] _T_52402; // @[Mux.scala 19:72:@25068.4]
  wire [15:0] _T_52404; // @[Mux.scala 19:72:@25069.4]
  wire [7:0] _T_52411; // @[Mux.scala 19:72:@25076.4]
  wire [7:0] _T_52418; // @[Mux.scala 19:72:@25083.4]
  wire [15:0] _T_52419; // @[Mux.scala 19:72:@25084.4]
  wire [15:0] _T_52421; // @[Mux.scala 19:72:@25085.4]
  wire [7:0] _T_52428; // @[Mux.scala 19:72:@25092.4]
  wire [7:0] _T_52435; // @[Mux.scala 19:72:@25099.4]
  wire [15:0] _T_52436; // @[Mux.scala 19:72:@25100.4]
  wire [15:0] _T_52438; // @[Mux.scala 19:72:@25101.4]
  wire [7:0] _T_52445; // @[Mux.scala 19:72:@25108.4]
  wire [7:0] _T_52452; // @[Mux.scala 19:72:@25115.4]
  wire [15:0] _T_52453; // @[Mux.scala 19:72:@25116.4]
  wire [15:0] _T_52455; // @[Mux.scala 19:72:@25117.4]
  wire [15:0] _T_52470; // @[Mux.scala 19:72:@25132.4]
  wire [15:0] _T_52472; // @[Mux.scala 19:72:@25133.4]
  wire [15:0] _T_52487; // @[Mux.scala 19:72:@25148.4]
  wire [15:0] _T_52489; // @[Mux.scala 19:72:@25149.4]
  wire [15:0] _T_52504; // @[Mux.scala 19:72:@25164.4]
  wire [15:0] _T_52506; // @[Mux.scala 19:72:@25165.4]
  wire [15:0] _T_52521; // @[Mux.scala 19:72:@25180.4]
  wire [15:0] _T_52523; // @[Mux.scala 19:72:@25181.4]
  wire [15:0] _T_52538; // @[Mux.scala 19:72:@25196.4]
  wire [15:0] _T_52540; // @[Mux.scala 19:72:@25197.4]
  wire [15:0] _T_52555; // @[Mux.scala 19:72:@25212.4]
  wire [15:0] _T_52557; // @[Mux.scala 19:72:@25213.4]
  wire [15:0] _T_52572; // @[Mux.scala 19:72:@25228.4]
  wire [15:0] _T_52574; // @[Mux.scala 19:72:@25229.4]
  wire [15:0] _T_52589; // @[Mux.scala 19:72:@25244.4]
  wire [15:0] _T_52591; // @[Mux.scala 19:72:@25245.4]
  wire [15:0] _T_52592; // @[Mux.scala 19:72:@25246.4]
  wire [15:0] _T_52593; // @[Mux.scala 19:72:@25247.4]
  wire [15:0] _T_52594; // @[Mux.scala 19:72:@25248.4]
  wire [15:0] _T_52595; // @[Mux.scala 19:72:@25249.4]
  wire [15:0] _T_52596; // @[Mux.scala 19:72:@25250.4]
  wire [15:0] _T_52597; // @[Mux.scala 19:72:@25251.4]
  wire [15:0] _T_52598; // @[Mux.scala 19:72:@25252.4]
  wire [15:0] _T_52599; // @[Mux.scala 19:72:@25253.4]
  wire [15:0] _T_52600; // @[Mux.scala 19:72:@25254.4]
  wire [15:0] _T_52601; // @[Mux.scala 19:72:@25255.4]
  wire [15:0] _T_52602; // @[Mux.scala 19:72:@25256.4]
  wire [15:0] _T_52603; // @[Mux.scala 19:72:@25257.4]
  wire [15:0] _T_52604; // @[Mux.scala 19:72:@25258.4]
  wire [15:0] _T_52605; // @[Mux.scala 19:72:@25259.4]
  wire [15:0] _T_52606; // @[Mux.scala 19:72:@25260.4]
  wire [7:0] _T_53184; // @[Mux.scala 19:72:@25610.4]
  wire [7:0] _T_53191; // @[Mux.scala 19:72:@25617.4]
  wire [15:0] _T_53192; // @[Mux.scala 19:72:@25618.4]
  wire [15:0] _T_53194; // @[Mux.scala 19:72:@25619.4]
  wire [7:0] _T_53201; // @[Mux.scala 19:72:@25626.4]
  wire [7:0] _T_53208; // @[Mux.scala 19:72:@25633.4]
  wire [15:0] _T_53209; // @[Mux.scala 19:72:@25634.4]
  wire [15:0] _T_53211; // @[Mux.scala 19:72:@25635.4]
  wire [7:0] _T_53218; // @[Mux.scala 19:72:@25642.4]
  wire [7:0] _T_53225; // @[Mux.scala 19:72:@25649.4]
  wire [15:0] _T_53226; // @[Mux.scala 19:72:@25650.4]
  wire [15:0] _T_53228; // @[Mux.scala 19:72:@25651.4]
  wire [7:0] _T_53235; // @[Mux.scala 19:72:@25658.4]
  wire [7:0] _T_53242; // @[Mux.scala 19:72:@25665.4]
  wire [15:0] _T_53243; // @[Mux.scala 19:72:@25666.4]
  wire [15:0] _T_53245; // @[Mux.scala 19:72:@25667.4]
  wire [7:0] _T_53252; // @[Mux.scala 19:72:@25674.4]
  wire [7:0] _T_53259; // @[Mux.scala 19:72:@25681.4]
  wire [15:0] _T_53260; // @[Mux.scala 19:72:@25682.4]
  wire [15:0] _T_53262; // @[Mux.scala 19:72:@25683.4]
  wire [7:0] _T_53269; // @[Mux.scala 19:72:@25690.4]
  wire [7:0] _T_53276; // @[Mux.scala 19:72:@25697.4]
  wire [15:0] _T_53277; // @[Mux.scala 19:72:@25698.4]
  wire [15:0] _T_53279; // @[Mux.scala 19:72:@25699.4]
  wire [7:0] _T_53286; // @[Mux.scala 19:72:@25706.4]
  wire [7:0] _T_53293; // @[Mux.scala 19:72:@25713.4]
  wire [15:0] _T_53294; // @[Mux.scala 19:72:@25714.4]
  wire [15:0] _T_53296; // @[Mux.scala 19:72:@25715.4]
  wire [7:0] _T_53303; // @[Mux.scala 19:72:@25722.4]
  wire [7:0] _T_53310; // @[Mux.scala 19:72:@25729.4]
  wire [15:0] _T_53311; // @[Mux.scala 19:72:@25730.4]
  wire [15:0] _T_53313; // @[Mux.scala 19:72:@25731.4]
  wire [15:0] _T_53328; // @[Mux.scala 19:72:@25746.4]
  wire [15:0] _T_53330; // @[Mux.scala 19:72:@25747.4]
  wire [15:0] _T_53345; // @[Mux.scala 19:72:@25762.4]
  wire [15:0] _T_53347; // @[Mux.scala 19:72:@25763.4]
  wire [15:0] _T_53362; // @[Mux.scala 19:72:@25778.4]
  wire [15:0] _T_53364; // @[Mux.scala 19:72:@25779.4]
  wire [15:0] _T_53379; // @[Mux.scala 19:72:@25794.4]
  wire [15:0] _T_53381; // @[Mux.scala 19:72:@25795.4]
  wire [15:0] _T_53396; // @[Mux.scala 19:72:@25810.4]
  wire [15:0] _T_53398; // @[Mux.scala 19:72:@25811.4]
  wire [15:0] _T_53413; // @[Mux.scala 19:72:@25826.4]
  wire [15:0] _T_53415; // @[Mux.scala 19:72:@25827.4]
  wire [15:0] _T_53430; // @[Mux.scala 19:72:@25842.4]
  wire [15:0] _T_53432; // @[Mux.scala 19:72:@25843.4]
  wire [15:0] _T_53447; // @[Mux.scala 19:72:@25858.4]
  wire [15:0] _T_53449; // @[Mux.scala 19:72:@25859.4]
  wire [15:0] _T_53450; // @[Mux.scala 19:72:@25860.4]
  wire [15:0] _T_53451; // @[Mux.scala 19:72:@25861.4]
  wire [15:0] _T_53452; // @[Mux.scala 19:72:@25862.4]
  wire [15:0] _T_53453; // @[Mux.scala 19:72:@25863.4]
  wire [15:0] _T_53454; // @[Mux.scala 19:72:@25864.4]
  wire [15:0] _T_53455; // @[Mux.scala 19:72:@25865.4]
  wire [15:0] _T_53456; // @[Mux.scala 19:72:@25866.4]
  wire [15:0] _T_53457; // @[Mux.scala 19:72:@25867.4]
  wire [15:0] _T_53458; // @[Mux.scala 19:72:@25868.4]
  wire [15:0] _T_53459; // @[Mux.scala 19:72:@25869.4]
  wire [15:0] _T_53460; // @[Mux.scala 19:72:@25870.4]
  wire [15:0] _T_53461; // @[Mux.scala 19:72:@25871.4]
  wire [15:0] _T_53462; // @[Mux.scala 19:72:@25872.4]
  wire [15:0] _T_53463; // @[Mux.scala 19:72:@25873.4]
  wire [15:0] _T_53464; // @[Mux.scala 19:72:@25874.4]
  wire [7:0] _T_54042; // @[Mux.scala 19:72:@26224.4]
  wire [7:0] _T_54049; // @[Mux.scala 19:72:@26231.4]
  wire [15:0] _T_54050; // @[Mux.scala 19:72:@26232.4]
  wire [15:0] _T_54052; // @[Mux.scala 19:72:@26233.4]
  wire [7:0] _T_54059; // @[Mux.scala 19:72:@26240.4]
  wire [7:0] _T_54066; // @[Mux.scala 19:72:@26247.4]
  wire [15:0] _T_54067; // @[Mux.scala 19:72:@26248.4]
  wire [15:0] _T_54069; // @[Mux.scala 19:72:@26249.4]
  wire [7:0] _T_54076; // @[Mux.scala 19:72:@26256.4]
  wire [7:0] _T_54083; // @[Mux.scala 19:72:@26263.4]
  wire [15:0] _T_54084; // @[Mux.scala 19:72:@26264.4]
  wire [15:0] _T_54086; // @[Mux.scala 19:72:@26265.4]
  wire [7:0] _T_54093; // @[Mux.scala 19:72:@26272.4]
  wire [7:0] _T_54100; // @[Mux.scala 19:72:@26279.4]
  wire [15:0] _T_54101; // @[Mux.scala 19:72:@26280.4]
  wire [15:0] _T_54103; // @[Mux.scala 19:72:@26281.4]
  wire [7:0] _T_54110; // @[Mux.scala 19:72:@26288.4]
  wire [7:0] _T_54117; // @[Mux.scala 19:72:@26295.4]
  wire [15:0] _T_54118; // @[Mux.scala 19:72:@26296.4]
  wire [15:0] _T_54120; // @[Mux.scala 19:72:@26297.4]
  wire [7:0] _T_54127; // @[Mux.scala 19:72:@26304.4]
  wire [7:0] _T_54134; // @[Mux.scala 19:72:@26311.4]
  wire [15:0] _T_54135; // @[Mux.scala 19:72:@26312.4]
  wire [15:0] _T_54137; // @[Mux.scala 19:72:@26313.4]
  wire [7:0] _T_54144; // @[Mux.scala 19:72:@26320.4]
  wire [7:0] _T_54151; // @[Mux.scala 19:72:@26327.4]
  wire [15:0] _T_54152; // @[Mux.scala 19:72:@26328.4]
  wire [15:0] _T_54154; // @[Mux.scala 19:72:@26329.4]
  wire [7:0] _T_54161; // @[Mux.scala 19:72:@26336.4]
  wire [7:0] _T_54168; // @[Mux.scala 19:72:@26343.4]
  wire [15:0] _T_54169; // @[Mux.scala 19:72:@26344.4]
  wire [15:0] _T_54171; // @[Mux.scala 19:72:@26345.4]
  wire [15:0] _T_54186; // @[Mux.scala 19:72:@26360.4]
  wire [15:0] _T_54188; // @[Mux.scala 19:72:@26361.4]
  wire [15:0] _T_54203; // @[Mux.scala 19:72:@26376.4]
  wire [15:0] _T_54205; // @[Mux.scala 19:72:@26377.4]
  wire [15:0] _T_54220; // @[Mux.scala 19:72:@26392.4]
  wire [15:0] _T_54222; // @[Mux.scala 19:72:@26393.4]
  wire [15:0] _T_54237; // @[Mux.scala 19:72:@26408.4]
  wire [15:0] _T_54239; // @[Mux.scala 19:72:@26409.4]
  wire [15:0] _T_54254; // @[Mux.scala 19:72:@26424.4]
  wire [15:0] _T_54256; // @[Mux.scala 19:72:@26425.4]
  wire [15:0] _T_54271; // @[Mux.scala 19:72:@26440.4]
  wire [15:0] _T_54273; // @[Mux.scala 19:72:@26441.4]
  wire [15:0] _T_54288; // @[Mux.scala 19:72:@26456.4]
  wire [15:0] _T_54290; // @[Mux.scala 19:72:@26457.4]
  wire [15:0] _T_54305; // @[Mux.scala 19:72:@26472.4]
  wire [15:0] _T_54307; // @[Mux.scala 19:72:@26473.4]
  wire [15:0] _T_54308; // @[Mux.scala 19:72:@26474.4]
  wire [15:0] _T_54309; // @[Mux.scala 19:72:@26475.4]
  wire [15:0] _T_54310; // @[Mux.scala 19:72:@26476.4]
  wire [15:0] _T_54311; // @[Mux.scala 19:72:@26477.4]
  wire [15:0] _T_54312; // @[Mux.scala 19:72:@26478.4]
  wire [15:0] _T_54313; // @[Mux.scala 19:72:@26479.4]
  wire [15:0] _T_54314; // @[Mux.scala 19:72:@26480.4]
  wire [15:0] _T_54315; // @[Mux.scala 19:72:@26481.4]
  wire [15:0] _T_54316; // @[Mux.scala 19:72:@26482.4]
  wire [15:0] _T_54317; // @[Mux.scala 19:72:@26483.4]
  wire [15:0] _T_54318; // @[Mux.scala 19:72:@26484.4]
  wire [15:0] _T_54319; // @[Mux.scala 19:72:@26485.4]
  wire [15:0] _T_54320; // @[Mux.scala 19:72:@26486.4]
  wire [15:0] _T_54321; // @[Mux.scala 19:72:@26487.4]
  wire [15:0] _T_54322; // @[Mux.scala 19:72:@26488.4]
  wire [7:0] _T_54900; // @[Mux.scala 19:72:@26838.4]
  wire [7:0] _T_54907; // @[Mux.scala 19:72:@26845.4]
  wire [15:0] _T_54908; // @[Mux.scala 19:72:@26846.4]
  wire [15:0] _T_54910; // @[Mux.scala 19:72:@26847.4]
  wire [7:0] _T_54917; // @[Mux.scala 19:72:@26854.4]
  wire [7:0] _T_54924; // @[Mux.scala 19:72:@26861.4]
  wire [15:0] _T_54925; // @[Mux.scala 19:72:@26862.4]
  wire [15:0] _T_54927; // @[Mux.scala 19:72:@26863.4]
  wire [7:0] _T_54934; // @[Mux.scala 19:72:@26870.4]
  wire [7:0] _T_54941; // @[Mux.scala 19:72:@26877.4]
  wire [15:0] _T_54942; // @[Mux.scala 19:72:@26878.4]
  wire [15:0] _T_54944; // @[Mux.scala 19:72:@26879.4]
  wire [7:0] _T_54951; // @[Mux.scala 19:72:@26886.4]
  wire [7:0] _T_54958; // @[Mux.scala 19:72:@26893.4]
  wire [15:0] _T_54959; // @[Mux.scala 19:72:@26894.4]
  wire [15:0] _T_54961; // @[Mux.scala 19:72:@26895.4]
  wire [7:0] _T_54968; // @[Mux.scala 19:72:@26902.4]
  wire [7:0] _T_54975; // @[Mux.scala 19:72:@26909.4]
  wire [15:0] _T_54976; // @[Mux.scala 19:72:@26910.4]
  wire [15:0] _T_54978; // @[Mux.scala 19:72:@26911.4]
  wire [7:0] _T_54985; // @[Mux.scala 19:72:@26918.4]
  wire [7:0] _T_54992; // @[Mux.scala 19:72:@26925.4]
  wire [15:0] _T_54993; // @[Mux.scala 19:72:@26926.4]
  wire [15:0] _T_54995; // @[Mux.scala 19:72:@26927.4]
  wire [7:0] _T_55002; // @[Mux.scala 19:72:@26934.4]
  wire [7:0] _T_55009; // @[Mux.scala 19:72:@26941.4]
  wire [15:0] _T_55010; // @[Mux.scala 19:72:@26942.4]
  wire [15:0] _T_55012; // @[Mux.scala 19:72:@26943.4]
  wire [7:0] _T_55019; // @[Mux.scala 19:72:@26950.4]
  wire [7:0] _T_55026; // @[Mux.scala 19:72:@26957.4]
  wire [15:0] _T_55027; // @[Mux.scala 19:72:@26958.4]
  wire [15:0] _T_55029; // @[Mux.scala 19:72:@26959.4]
  wire [15:0] _T_55044; // @[Mux.scala 19:72:@26974.4]
  wire [15:0] _T_55046; // @[Mux.scala 19:72:@26975.4]
  wire [15:0] _T_55061; // @[Mux.scala 19:72:@26990.4]
  wire [15:0] _T_55063; // @[Mux.scala 19:72:@26991.4]
  wire [15:0] _T_55078; // @[Mux.scala 19:72:@27006.4]
  wire [15:0] _T_55080; // @[Mux.scala 19:72:@27007.4]
  wire [15:0] _T_55095; // @[Mux.scala 19:72:@27022.4]
  wire [15:0] _T_55097; // @[Mux.scala 19:72:@27023.4]
  wire [15:0] _T_55112; // @[Mux.scala 19:72:@27038.4]
  wire [15:0] _T_55114; // @[Mux.scala 19:72:@27039.4]
  wire [15:0] _T_55129; // @[Mux.scala 19:72:@27054.4]
  wire [15:0] _T_55131; // @[Mux.scala 19:72:@27055.4]
  wire [15:0] _T_55146; // @[Mux.scala 19:72:@27070.4]
  wire [15:0] _T_55148; // @[Mux.scala 19:72:@27071.4]
  wire [15:0] _T_55163; // @[Mux.scala 19:72:@27086.4]
  wire [15:0] _T_55165; // @[Mux.scala 19:72:@27087.4]
  wire [15:0] _T_55166; // @[Mux.scala 19:72:@27088.4]
  wire [15:0] _T_55167; // @[Mux.scala 19:72:@27089.4]
  wire [15:0] _T_55168; // @[Mux.scala 19:72:@27090.4]
  wire [15:0] _T_55169; // @[Mux.scala 19:72:@27091.4]
  wire [15:0] _T_55170; // @[Mux.scala 19:72:@27092.4]
  wire [15:0] _T_55171; // @[Mux.scala 19:72:@27093.4]
  wire [15:0] _T_55172; // @[Mux.scala 19:72:@27094.4]
  wire [15:0] _T_55173; // @[Mux.scala 19:72:@27095.4]
  wire [15:0] _T_55174; // @[Mux.scala 19:72:@27096.4]
  wire [15:0] _T_55175; // @[Mux.scala 19:72:@27097.4]
  wire [15:0] _T_55176; // @[Mux.scala 19:72:@27098.4]
  wire [15:0] _T_55177; // @[Mux.scala 19:72:@27099.4]
  wire [15:0] _T_55178; // @[Mux.scala 19:72:@27100.4]
  wire [15:0] _T_55179; // @[Mux.scala 19:72:@27101.4]
  wire [15:0] _T_55180; // @[Mux.scala 19:72:@27102.4]
  wire [7:0] _T_55758; // @[Mux.scala 19:72:@27452.4]
  wire [7:0] _T_55765; // @[Mux.scala 19:72:@27459.4]
  wire [15:0] _T_55766; // @[Mux.scala 19:72:@27460.4]
  wire [15:0] _T_55768; // @[Mux.scala 19:72:@27461.4]
  wire [7:0] _T_55775; // @[Mux.scala 19:72:@27468.4]
  wire [7:0] _T_55782; // @[Mux.scala 19:72:@27475.4]
  wire [15:0] _T_55783; // @[Mux.scala 19:72:@27476.4]
  wire [15:0] _T_55785; // @[Mux.scala 19:72:@27477.4]
  wire [7:0] _T_55792; // @[Mux.scala 19:72:@27484.4]
  wire [7:0] _T_55799; // @[Mux.scala 19:72:@27491.4]
  wire [15:0] _T_55800; // @[Mux.scala 19:72:@27492.4]
  wire [15:0] _T_55802; // @[Mux.scala 19:72:@27493.4]
  wire [7:0] _T_55809; // @[Mux.scala 19:72:@27500.4]
  wire [7:0] _T_55816; // @[Mux.scala 19:72:@27507.4]
  wire [15:0] _T_55817; // @[Mux.scala 19:72:@27508.4]
  wire [15:0] _T_55819; // @[Mux.scala 19:72:@27509.4]
  wire [7:0] _T_55826; // @[Mux.scala 19:72:@27516.4]
  wire [7:0] _T_55833; // @[Mux.scala 19:72:@27523.4]
  wire [15:0] _T_55834; // @[Mux.scala 19:72:@27524.4]
  wire [15:0] _T_55836; // @[Mux.scala 19:72:@27525.4]
  wire [7:0] _T_55843; // @[Mux.scala 19:72:@27532.4]
  wire [7:0] _T_55850; // @[Mux.scala 19:72:@27539.4]
  wire [15:0] _T_55851; // @[Mux.scala 19:72:@27540.4]
  wire [15:0] _T_55853; // @[Mux.scala 19:72:@27541.4]
  wire [7:0] _T_55860; // @[Mux.scala 19:72:@27548.4]
  wire [7:0] _T_55867; // @[Mux.scala 19:72:@27555.4]
  wire [15:0] _T_55868; // @[Mux.scala 19:72:@27556.4]
  wire [15:0] _T_55870; // @[Mux.scala 19:72:@27557.4]
  wire [7:0] _T_55877; // @[Mux.scala 19:72:@27564.4]
  wire [7:0] _T_55884; // @[Mux.scala 19:72:@27571.4]
  wire [15:0] _T_55885; // @[Mux.scala 19:72:@27572.4]
  wire [15:0] _T_55887; // @[Mux.scala 19:72:@27573.4]
  wire [15:0] _T_55902; // @[Mux.scala 19:72:@27588.4]
  wire [15:0] _T_55904; // @[Mux.scala 19:72:@27589.4]
  wire [15:0] _T_55919; // @[Mux.scala 19:72:@27604.4]
  wire [15:0] _T_55921; // @[Mux.scala 19:72:@27605.4]
  wire [15:0] _T_55936; // @[Mux.scala 19:72:@27620.4]
  wire [15:0] _T_55938; // @[Mux.scala 19:72:@27621.4]
  wire [15:0] _T_55953; // @[Mux.scala 19:72:@27636.4]
  wire [15:0] _T_55955; // @[Mux.scala 19:72:@27637.4]
  wire [15:0] _T_55970; // @[Mux.scala 19:72:@27652.4]
  wire [15:0] _T_55972; // @[Mux.scala 19:72:@27653.4]
  wire [15:0] _T_55987; // @[Mux.scala 19:72:@27668.4]
  wire [15:0] _T_55989; // @[Mux.scala 19:72:@27669.4]
  wire [15:0] _T_56004; // @[Mux.scala 19:72:@27684.4]
  wire [15:0] _T_56006; // @[Mux.scala 19:72:@27685.4]
  wire [15:0] _T_56021; // @[Mux.scala 19:72:@27700.4]
  wire [15:0] _T_56023; // @[Mux.scala 19:72:@27701.4]
  wire [15:0] _T_56024; // @[Mux.scala 19:72:@27702.4]
  wire [15:0] _T_56025; // @[Mux.scala 19:72:@27703.4]
  wire [15:0] _T_56026; // @[Mux.scala 19:72:@27704.4]
  wire [15:0] _T_56027; // @[Mux.scala 19:72:@27705.4]
  wire [15:0] _T_56028; // @[Mux.scala 19:72:@27706.4]
  wire [15:0] _T_56029; // @[Mux.scala 19:72:@27707.4]
  wire [15:0] _T_56030; // @[Mux.scala 19:72:@27708.4]
  wire [15:0] _T_56031; // @[Mux.scala 19:72:@27709.4]
  wire [15:0] _T_56032; // @[Mux.scala 19:72:@27710.4]
  wire [15:0] _T_56033; // @[Mux.scala 19:72:@27711.4]
  wire [15:0] _T_56034; // @[Mux.scala 19:72:@27712.4]
  wire [15:0] _T_56035; // @[Mux.scala 19:72:@27713.4]
  wire [15:0] _T_56036; // @[Mux.scala 19:72:@27714.4]
  wire [15:0] _T_56037; // @[Mux.scala 19:72:@27715.4]
  wire [15:0] _T_56038; // @[Mux.scala 19:72:@27716.4]
  wire [7:0] _T_56616; // @[Mux.scala 19:72:@28066.4]
  wire [7:0] _T_56623; // @[Mux.scala 19:72:@28073.4]
  wire [15:0] _T_56624; // @[Mux.scala 19:72:@28074.4]
  wire [15:0] _T_56626; // @[Mux.scala 19:72:@28075.4]
  wire [7:0] _T_56633; // @[Mux.scala 19:72:@28082.4]
  wire [7:0] _T_56640; // @[Mux.scala 19:72:@28089.4]
  wire [15:0] _T_56641; // @[Mux.scala 19:72:@28090.4]
  wire [15:0] _T_56643; // @[Mux.scala 19:72:@28091.4]
  wire [7:0] _T_56650; // @[Mux.scala 19:72:@28098.4]
  wire [7:0] _T_56657; // @[Mux.scala 19:72:@28105.4]
  wire [15:0] _T_56658; // @[Mux.scala 19:72:@28106.4]
  wire [15:0] _T_56660; // @[Mux.scala 19:72:@28107.4]
  wire [7:0] _T_56667; // @[Mux.scala 19:72:@28114.4]
  wire [7:0] _T_56674; // @[Mux.scala 19:72:@28121.4]
  wire [15:0] _T_56675; // @[Mux.scala 19:72:@28122.4]
  wire [15:0] _T_56677; // @[Mux.scala 19:72:@28123.4]
  wire [7:0] _T_56684; // @[Mux.scala 19:72:@28130.4]
  wire [7:0] _T_56691; // @[Mux.scala 19:72:@28137.4]
  wire [15:0] _T_56692; // @[Mux.scala 19:72:@28138.4]
  wire [15:0] _T_56694; // @[Mux.scala 19:72:@28139.4]
  wire [7:0] _T_56701; // @[Mux.scala 19:72:@28146.4]
  wire [7:0] _T_56708; // @[Mux.scala 19:72:@28153.4]
  wire [15:0] _T_56709; // @[Mux.scala 19:72:@28154.4]
  wire [15:0] _T_56711; // @[Mux.scala 19:72:@28155.4]
  wire [7:0] _T_56718; // @[Mux.scala 19:72:@28162.4]
  wire [7:0] _T_56725; // @[Mux.scala 19:72:@28169.4]
  wire [15:0] _T_56726; // @[Mux.scala 19:72:@28170.4]
  wire [15:0] _T_56728; // @[Mux.scala 19:72:@28171.4]
  wire [7:0] _T_56735; // @[Mux.scala 19:72:@28178.4]
  wire [7:0] _T_56742; // @[Mux.scala 19:72:@28185.4]
  wire [15:0] _T_56743; // @[Mux.scala 19:72:@28186.4]
  wire [15:0] _T_56745; // @[Mux.scala 19:72:@28187.4]
  wire [15:0] _T_56760; // @[Mux.scala 19:72:@28202.4]
  wire [15:0] _T_56762; // @[Mux.scala 19:72:@28203.4]
  wire [15:0] _T_56777; // @[Mux.scala 19:72:@28218.4]
  wire [15:0] _T_56779; // @[Mux.scala 19:72:@28219.4]
  wire [15:0] _T_56794; // @[Mux.scala 19:72:@28234.4]
  wire [15:0] _T_56796; // @[Mux.scala 19:72:@28235.4]
  wire [15:0] _T_56811; // @[Mux.scala 19:72:@28250.4]
  wire [15:0] _T_56813; // @[Mux.scala 19:72:@28251.4]
  wire [15:0] _T_56828; // @[Mux.scala 19:72:@28266.4]
  wire [15:0] _T_56830; // @[Mux.scala 19:72:@28267.4]
  wire [15:0] _T_56845; // @[Mux.scala 19:72:@28282.4]
  wire [15:0] _T_56847; // @[Mux.scala 19:72:@28283.4]
  wire [15:0] _T_56862; // @[Mux.scala 19:72:@28298.4]
  wire [15:0] _T_56864; // @[Mux.scala 19:72:@28299.4]
  wire [15:0] _T_56879; // @[Mux.scala 19:72:@28314.4]
  wire [15:0] _T_56881; // @[Mux.scala 19:72:@28315.4]
  wire [15:0] _T_56882; // @[Mux.scala 19:72:@28316.4]
  wire [15:0] _T_56883; // @[Mux.scala 19:72:@28317.4]
  wire [15:0] _T_56884; // @[Mux.scala 19:72:@28318.4]
  wire [15:0] _T_56885; // @[Mux.scala 19:72:@28319.4]
  wire [15:0] _T_56886; // @[Mux.scala 19:72:@28320.4]
  wire [15:0] _T_56887; // @[Mux.scala 19:72:@28321.4]
  wire [15:0] _T_56888; // @[Mux.scala 19:72:@28322.4]
  wire [15:0] _T_56889; // @[Mux.scala 19:72:@28323.4]
  wire [15:0] _T_56890; // @[Mux.scala 19:72:@28324.4]
  wire [15:0] _T_56891; // @[Mux.scala 19:72:@28325.4]
  wire [15:0] _T_56892; // @[Mux.scala 19:72:@28326.4]
  wire [15:0] _T_56893; // @[Mux.scala 19:72:@28327.4]
  wire [15:0] _T_56894; // @[Mux.scala 19:72:@28328.4]
  wire [15:0] _T_56895; // @[Mux.scala 19:72:@28329.4]
  wire [15:0] _T_56896; // @[Mux.scala 19:72:@28330.4]
  wire [7:0] _T_57474; // @[Mux.scala 19:72:@28680.4]
  wire [7:0] _T_57481; // @[Mux.scala 19:72:@28687.4]
  wire [15:0] _T_57482; // @[Mux.scala 19:72:@28688.4]
  wire [15:0] _T_57484; // @[Mux.scala 19:72:@28689.4]
  wire [7:0] _T_57491; // @[Mux.scala 19:72:@28696.4]
  wire [7:0] _T_57498; // @[Mux.scala 19:72:@28703.4]
  wire [15:0] _T_57499; // @[Mux.scala 19:72:@28704.4]
  wire [15:0] _T_57501; // @[Mux.scala 19:72:@28705.4]
  wire [7:0] _T_57508; // @[Mux.scala 19:72:@28712.4]
  wire [7:0] _T_57515; // @[Mux.scala 19:72:@28719.4]
  wire [15:0] _T_57516; // @[Mux.scala 19:72:@28720.4]
  wire [15:0] _T_57518; // @[Mux.scala 19:72:@28721.4]
  wire [7:0] _T_57525; // @[Mux.scala 19:72:@28728.4]
  wire [7:0] _T_57532; // @[Mux.scala 19:72:@28735.4]
  wire [15:0] _T_57533; // @[Mux.scala 19:72:@28736.4]
  wire [15:0] _T_57535; // @[Mux.scala 19:72:@28737.4]
  wire [7:0] _T_57542; // @[Mux.scala 19:72:@28744.4]
  wire [7:0] _T_57549; // @[Mux.scala 19:72:@28751.4]
  wire [15:0] _T_57550; // @[Mux.scala 19:72:@28752.4]
  wire [15:0] _T_57552; // @[Mux.scala 19:72:@28753.4]
  wire [7:0] _T_57559; // @[Mux.scala 19:72:@28760.4]
  wire [7:0] _T_57566; // @[Mux.scala 19:72:@28767.4]
  wire [15:0] _T_57567; // @[Mux.scala 19:72:@28768.4]
  wire [15:0] _T_57569; // @[Mux.scala 19:72:@28769.4]
  wire [7:0] _T_57576; // @[Mux.scala 19:72:@28776.4]
  wire [7:0] _T_57583; // @[Mux.scala 19:72:@28783.4]
  wire [15:0] _T_57584; // @[Mux.scala 19:72:@28784.4]
  wire [15:0] _T_57586; // @[Mux.scala 19:72:@28785.4]
  wire [7:0] _T_57593; // @[Mux.scala 19:72:@28792.4]
  wire [7:0] _T_57600; // @[Mux.scala 19:72:@28799.4]
  wire [15:0] _T_57601; // @[Mux.scala 19:72:@28800.4]
  wire [15:0] _T_57603; // @[Mux.scala 19:72:@28801.4]
  wire [15:0] _T_57618; // @[Mux.scala 19:72:@28816.4]
  wire [15:0] _T_57620; // @[Mux.scala 19:72:@28817.4]
  wire [15:0] _T_57635; // @[Mux.scala 19:72:@28832.4]
  wire [15:0] _T_57637; // @[Mux.scala 19:72:@28833.4]
  wire [15:0] _T_57652; // @[Mux.scala 19:72:@28848.4]
  wire [15:0] _T_57654; // @[Mux.scala 19:72:@28849.4]
  wire [15:0] _T_57669; // @[Mux.scala 19:72:@28864.4]
  wire [15:0] _T_57671; // @[Mux.scala 19:72:@28865.4]
  wire [15:0] _T_57686; // @[Mux.scala 19:72:@28880.4]
  wire [15:0] _T_57688; // @[Mux.scala 19:72:@28881.4]
  wire [15:0] _T_57703; // @[Mux.scala 19:72:@28896.4]
  wire [15:0] _T_57705; // @[Mux.scala 19:72:@28897.4]
  wire [15:0] _T_57720; // @[Mux.scala 19:72:@28912.4]
  wire [15:0] _T_57722; // @[Mux.scala 19:72:@28913.4]
  wire [15:0] _T_57737; // @[Mux.scala 19:72:@28928.4]
  wire [15:0] _T_57739; // @[Mux.scala 19:72:@28929.4]
  wire [15:0] _T_57740; // @[Mux.scala 19:72:@28930.4]
  wire [15:0] _T_57741; // @[Mux.scala 19:72:@28931.4]
  wire [15:0] _T_57742; // @[Mux.scala 19:72:@28932.4]
  wire [15:0] _T_57743; // @[Mux.scala 19:72:@28933.4]
  wire [15:0] _T_57744; // @[Mux.scala 19:72:@28934.4]
  wire [15:0] _T_57745; // @[Mux.scala 19:72:@28935.4]
  wire [15:0] _T_57746; // @[Mux.scala 19:72:@28936.4]
  wire [15:0] _T_57747; // @[Mux.scala 19:72:@28937.4]
  wire [15:0] _T_57748; // @[Mux.scala 19:72:@28938.4]
  wire [15:0] _T_57749; // @[Mux.scala 19:72:@28939.4]
  wire [15:0] _T_57750; // @[Mux.scala 19:72:@28940.4]
  wire [15:0] _T_57751; // @[Mux.scala 19:72:@28941.4]
  wire [15:0] _T_57752; // @[Mux.scala 19:72:@28942.4]
  wire [15:0] _T_57753; // @[Mux.scala 19:72:@28943.4]
  wire [15:0] _T_57754; // @[Mux.scala 19:72:@28944.4]
  wire [7:0] _T_58332; // @[Mux.scala 19:72:@29294.4]
  wire [7:0] _T_58339; // @[Mux.scala 19:72:@29301.4]
  wire [15:0] _T_58340; // @[Mux.scala 19:72:@29302.4]
  wire [15:0] _T_58342; // @[Mux.scala 19:72:@29303.4]
  wire [7:0] _T_58349; // @[Mux.scala 19:72:@29310.4]
  wire [7:0] _T_58356; // @[Mux.scala 19:72:@29317.4]
  wire [15:0] _T_58357; // @[Mux.scala 19:72:@29318.4]
  wire [15:0] _T_58359; // @[Mux.scala 19:72:@29319.4]
  wire [7:0] _T_58366; // @[Mux.scala 19:72:@29326.4]
  wire [7:0] _T_58373; // @[Mux.scala 19:72:@29333.4]
  wire [15:0] _T_58374; // @[Mux.scala 19:72:@29334.4]
  wire [15:0] _T_58376; // @[Mux.scala 19:72:@29335.4]
  wire [7:0] _T_58383; // @[Mux.scala 19:72:@29342.4]
  wire [7:0] _T_58390; // @[Mux.scala 19:72:@29349.4]
  wire [15:0] _T_58391; // @[Mux.scala 19:72:@29350.4]
  wire [15:0] _T_58393; // @[Mux.scala 19:72:@29351.4]
  wire [7:0] _T_58400; // @[Mux.scala 19:72:@29358.4]
  wire [7:0] _T_58407; // @[Mux.scala 19:72:@29365.4]
  wire [15:0] _T_58408; // @[Mux.scala 19:72:@29366.4]
  wire [15:0] _T_58410; // @[Mux.scala 19:72:@29367.4]
  wire [7:0] _T_58417; // @[Mux.scala 19:72:@29374.4]
  wire [7:0] _T_58424; // @[Mux.scala 19:72:@29381.4]
  wire [15:0] _T_58425; // @[Mux.scala 19:72:@29382.4]
  wire [15:0] _T_58427; // @[Mux.scala 19:72:@29383.4]
  wire [7:0] _T_58434; // @[Mux.scala 19:72:@29390.4]
  wire [7:0] _T_58441; // @[Mux.scala 19:72:@29397.4]
  wire [15:0] _T_58442; // @[Mux.scala 19:72:@29398.4]
  wire [15:0] _T_58444; // @[Mux.scala 19:72:@29399.4]
  wire [7:0] _T_58451; // @[Mux.scala 19:72:@29406.4]
  wire [7:0] _T_58458; // @[Mux.scala 19:72:@29413.4]
  wire [15:0] _T_58459; // @[Mux.scala 19:72:@29414.4]
  wire [15:0] _T_58461; // @[Mux.scala 19:72:@29415.4]
  wire [15:0] _T_58476; // @[Mux.scala 19:72:@29430.4]
  wire [15:0] _T_58478; // @[Mux.scala 19:72:@29431.4]
  wire [15:0] _T_58493; // @[Mux.scala 19:72:@29446.4]
  wire [15:0] _T_58495; // @[Mux.scala 19:72:@29447.4]
  wire [15:0] _T_58510; // @[Mux.scala 19:72:@29462.4]
  wire [15:0] _T_58512; // @[Mux.scala 19:72:@29463.4]
  wire [15:0] _T_58527; // @[Mux.scala 19:72:@29478.4]
  wire [15:0] _T_58529; // @[Mux.scala 19:72:@29479.4]
  wire [15:0] _T_58544; // @[Mux.scala 19:72:@29494.4]
  wire [15:0] _T_58546; // @[Mux.scala 19:72:@29495.4]
  wire [15:0] _T_58561; // @[Mux.scala 19:72:@29510.4]
  wire [15:0] _T_58563; // @[Mux.scala 19:72:@29511.4]
  wire [15:0] _T_58578; // @[Mux.scala 19:72:@29526.4]
  wire [15:0] _T_58580; // @[Mux.scala 19:72:@29527.4]
  wire [15:0] _T_58595; // @[Mux.scala 19:72:@29542.4]
  wire [15:0] _T_58597; // @[Mux.scala 19:72:@29543.4]
  wire [15:0] _T_58598; // @[Mux.scala 19:72:@29544.4]
  wire [15:0] _T_58599; // @[Mux.scala 19:72:@29545.4]
  wire [15:0] _T_58600; // @[Mux.scala 19:72:@29546.4]
  wire [15:0] _T_58601; // @[Mux.scala 19:72:@29547.4]
  wire [15:0] _T_58602; // @[Mux.scala 19:72:@29548.4]
  wire [15:0] _T_58603; // @[Mux.scala 19:72:@29549.4]
  wire [15:0] _T_58604; // @[Mux.scala 19:72:@29550.4]
  wire [15:0] _T_58605; // @[Mux.scala 19:72:@29551.4]
  wire [15:0] _T_58606; // @[Mux.scala 19:72:@29552.4]
  wire [15:0] _T_58607; // @[Mux.scala 19:72:@29553.4]
  wire [15:0] _T_58608; // @[Mux.scala 19:72:@29554.4]
  wire [15:0] _T_58609; // @[Mux.scala 19:72:@29555.4]
  wire [15:0] _T_58610; // @[Mux.scala 19:72:@29556.4]
  wire [15:0] _T_58611; // @[Mux.scala 19:72:@29557.4]
  wire [15:0] _T_58612; // @[Mux.scala 19:72:@29558.4]
  wire [7:0] _T_59190; // @[Mux.scala 19:72:@29908.4]
  wire [7:0] _T_59197; // @[Mux.scala 19:72:@29915.4]
  wire [15:0] _T_59198; // @[Mux.scala 19:72:@29916.4]
  wire [15:0] _T_59200; // @[Mux.scala 19:72:@29917.4]
  wire [7:0] _T_59207; // @[Mux.scala 19:72:@29924.4]
  wire [7:0] _T_59214; // @[Mux.scala 19:72:@29931.4]
  wire [15:0] _T_59215; // @[Mux.scala 19:72:@29932.4]
  wire [15:0] _T_59217; // @[Mux.scala 19:72:@29933.4]
  wire [7:0] _T_59224; // @[Mux.scala 19:72:@29940.4]
  wire [7:0] _T_59231; // @[Mux.scala 19:72:@29947.4]
  wire [15:0] _T_59232; // @[Mux.scala 19:72:@29948.4]
  wire [15:0] _T_59234; // @[Mux.scala 19:72:@29949.4]
  wire [7:0] _T_59241; // @[Mux.scala 19:72:@29956.4]
  wire [7:0] _T_59248; // @[Mux.scala 19:72:@29963.4]
  wire [15:0] _T_59249; // @[Mux.scala 19:72:@29964.4]
  wire [15:0] _T_59251; // @[Mux.scala 19:72:@29965.4]
  wire [7:0] _T_59258; // @[Mux.scala 19:72:@29972.4]
  wire [7:0] _T_59265; // @[Mux.scala 19:72:@29979.4]
  wire [15:0] _T_59266; // @[Mux.scala 19:72:@29980.4]
  wire [15:0] _T_59268; // @[Mux.scala 19:72:@29981.4]
  wire [7:0] _T_59275; // @[Mux.scala 19:72:@29988.4]
  wire [7:0] _T_59282; // @[Mux.scala 19:72:@29995.4]
  wire [15:0] _T_59283; // @[Mux.scala 19:72:@29996.4]
  wire [15:0] _T_59285; // @[Mux.scala 19:72:@29997.4]
  wire [7:0] _T_59292; // @[Mux.scala 19:72:@30004.4]
  wire [7:0] _T_59299; // @[Mux.scala 19:72:@30011.4]
  wire [15:0] _T_59300; // @[Mux.scala 19:72:@30012.4]
  wire [15:0] _T_59302; // @[Mux.scala 19:72:@30013.4]
  wire [7:0] _T_59309; // @[Mux.scala 19:72:@30020.4]
  wire [7:0] _T_59316; // @[Mux.scala 19:72:@30027.4]
  wire [15:0] _T_59317; // @[Mux.scala 19:72:@30028.4]
  wire [15:0] _T_59319; // @[Mux.scala 19:72:@30029.4]
  wire [15:0] _T_59334; // @[Mux.scala 19:72:@30044.4]
  wire [15:0] _T_59336; // @[Mux.scala 19:72:@30045.4]
  wire [15:0] _T_59351; // @[Mux.scala 19:72:@30060.4]
  wire [15:0] _T_59353; // @[Mux.scala 19:72:@30061.4]
  wire [15:0] _T_59368; // @[Mux.scala 19:72:@30076.4]
  wire [15:0] _T_59370; // @[Mux.scala 19:72:@30077.4]
  wire [15:0] _T_59385; // @[Mux.scala 19:72:@30092.4]
  wire [15:0] _T_59387; // @[Mux.scala 19:72:@30093.4]
  wire [15:0] _T_59402; // @[Mux.scala 19:72:@30108.4]
  wire [15:0] _T_59404; // @[Mux.scala 19:72:@30109.4]
  wire [15:0] _T_59419; // @[Mux.scala 19:72:@30124.4]
  wire [15:0] _T_59421; // @[Mux.scala 19:72:@30125.4]
  wire [15:0] _T_59436; // @[Mux.scala 19:72:@30140.4]
  wire [15:0] _T_59438; // @[Mux.scala 19:72:@30141.4]
  wire [15:0] _T_59453; // @[Mux.scala 19:72:@30156.4]
  wire [15:0] _T_59455; // @[Mux.scala 19:72:@30157.4]
  wire [15:0] _T_59456; // @[Mux.scala 19:72:@30158.4]
  wire [15:0] _T_59457; // @[Mux.scala 19:72:@30159.4]
  wire [15:0] _T_59458; // @[Mux.scala 19:72:@30160.4]
  wire [15:0] _T_59459; // @[Mux.scala 19:72:@30161.4]
  wire [15:0] _T_59460; // @[Mux.scala 19:72:@30162.4]
  wire [15:0] _T_59461; // @[Mux.scala 19:72:@30163.4]
  wire [15:0] _T_59462; // @[Mux.scala 19:72:@30164.4]
  wire [15:0] _T_59463; // @[Mux.scala 19:72:@30165.4]
  wire [15:0] _T_59464; // @[Mux.scala 19:72:@30166.4]
  wire [15:0] _T_59465; // @[Mux.scala 19:72:@30167.4]
  wire [15:0] _T_59466; // @[Mux.scala 19:72:@30168.4]
  wire [15:0] _T_59467; // @[Mux.scala 19:72:@30169.4]
  wire [15:0] _T_59468; // @[Mux.scala 19:72:@30170.4]
  wire [15:0] _T_59469; // @[Mux.scala 19:72:@30171.4]
  wire [15:0] _T_59470; // @[Mux.scala 19:72:@30172.4]
  wire [7:0] _T_60048; // @[Mux.scala 19:72:@30522.4]
  wire [7:0] _T_60055; // @[Mux.scala 19:72:@30529.4]
  wire [15:0] _T_60056; // @[Mux.scala 19:72:@30530.4]
  wire [15:0] _T_60058; // @[Mux.scala 19:72:@30531.4]
  wire [7:0] _T_60065; // @[Mux.scala 19:72:@30538.4]
  wire [7:0] _T_60072; // @[Mux.scala 19:72:@30545.4]
  wire [15:0] _T_60073; // @[Mux.scala 19:72:@30546.4]
  wire [15:0] _T_60075; // @[Mux.scala 19:72:@30547.4]
  wire [7:0] _T_60082; // @[Mux.scala 19:72:@30554.4]
  wire [7:0] _T_60089; // @[Mux.scala 19:72:@30561.4]
  wire [15:0] _T_60090; // @[Mux.scala 19:72:@30562.4]
  wire [15:0] _T_60092; // @[Mux.scala 19:72:@30563.4]
  wire [7:0] _T_60099; // @[Mux.scala 19:72:@30570.4]
  wire [7:0] _T_60106; // @[Mux.scala 19:72:@30577.4]
  wire [15:0] _T_60107; // @[Mux.scala 19:72:@30578.4]
  wire [15:0] _T_60109; // @[Mux.scala 19:72:@30579.4]
  wire [7:0] _T_60116; // @[Mux.scala 19:72:@30586.4]
  wire [7:0] _T_60123; // @[Mux.scala 19:72:@30593.4]
  wire [15:0] _T_60124; // @[Mux.scala 19:72:@30594.4]
  wire [15:0] _T_60126; // @[Mux.scala 19:72:@30595.4]
  wire [7:0] _T_60133; // @[Mux.scala 19:72:@30602.4]
  wire [7:0] _T_60140; // @[Mux.scala 19:72:@30609.4]
  wire [15:0] _T_60141; // @[Mux.scala 19:72:@30610.4]
  wire [15:0] _T_60143; // @[Mux.scala 19:72:@30611.4]
  wire [7:0] _T_60150; // @[Mux.scala 19:72:@30618.4]
  wire [7:0] _T_60157; // @[Mux.scala 19:72:@30625.4]
  wire [15:0] _T_60158; // @[Mux.scala 19:72:@30626.4]
  wire [15:0] _T_60160; // @[Mux.scala 19:72:@30627.4]
  wire [7:0] _T_60167; // @[Mux.scala 19:72:@30634.4]
  wire [7:0] _T_60174; // @[Mux.scala 19:72:@30641.4]
  wire [15:0] _T_60175; // @[Mux.scala 19:72:@30642.4]
  wire [15:0] _T_60177; // @[Mux.scala 19:72:@30643.4]
  wire [15:0] _T_60192; // @[Mux.scala 19:72:@30658.4]
  wire [15:0] _T_60194; // @[Mux.scala 19:72:@30659.4]
  wire [15:0] _T_60209; // @[Mux.scala 19:72:@30674.4]
  wire [15:0] _T_60211; // @[Mux.scala 19:72:@30675.4]
  wire [15:0] _T_60226; // @[Mux.scala 19:72:@30690.4]
  wire [15:0] _T_60228; // @[Mux.scala 19:72:@30691.4]
  wire [15:0] _T_60243; // @[Mux.scala 19:72:@30706.4]
  wire [15:0] _T_60245; // @[Mux.scala 19:72:@30707.4]
  wire [15:0] _T_60260; // @[Mux.scala 19:72:@30722.4]
  wire [15:0] _T_60262; // @[Mux.scala 19:72:@30723.4]
  wire [15:0] _T_60277; // @[Mux.scala 19:72:@30738.4]
  wire [15:0] _T_60279; // @[Mux.scala 19:72:@30739.4]
  wire [15:0] _T_60294; // @[Mux.scala 19:72:@30754.4]
  wire [15:0] _T_60296; // @[Mux.scala 19:72:@30755.4]
  wire [15:0] _T_60311; // @[Mux.scala 19:72:@30770.4]
  wire [15:0] _T_60313; // @[Mux.scala 19:72:@30771.4]
  wire [15:0] _T_60314; // @[Mux.scala 19:72:@30772.4]
  wire [15:0] _T_60315; // @[Mux.scala 19:72:@30773.4]
  wire [15:0] _T_60316; // @[Mux.scala 19:72:@30774.4]
  wire [15:0] _T_60317; // @[Mux.scala 19:72:@30775.4]
  wire [15:0] _T_60318; // @[Mux.scala 19:72:@30776.4]
  wire [15:0] _T_60319; // @[Mux.scala 19:72:@30777.4]
  wire [15:0] _T_60320; // @[Mux.scala 19:72:@30778.4]
  wire [15:0] _T_60321; // @[Mux.scala 19:72:@30779.4]
  wire [15:0] _T_60322; // @[Mux.scala 19:72:@30780.4]
  wire [15:0] _T_60323; // @[Mux.scala 19:72:@30781.4]
  wire [15:0] _T_60324; // @[Mux.scala 19:72:@30782.4]
  wire [15:0] _T_60325; // @[Mux.scala 19:72:@30783.4]
  wire [15:0] _T_60326; // @[Mux.scala 19:72:@30784.4]
  wire [15:0] _T_60327; // @[Mux.scala 19:72:@30785.4]
  wire [15:0] _T_60328; // @[Mux.scala 19:72:@30786.4]
  wire [7:0] _T_60906; // @[Mux.scala 19:72:@31136.4]
  wire [7:0] _T_60913; // @[Mux.scala 19:72:@31143.4]
  wire [15:0] _T_60914; // @[Mux.scala 19:72:@31144.4]
  wire [15:0] _T_60916; // @[Mux.scala 19:72:@31145.4]
  wire [7:0] _T_60923; // @[Mux.scala 19:72:@31152.4]
  wire [7:0] _T_60930; // @[Mux.scala 19:72:@31159.4]
  wire [15:0] _T_60931; // @[Mux.scala 19:72:@31160.4]
  wire [15:0] _T_60933; // @[Mux.scala 19:72:@31161.4]
  wire [7:0] _T_60940; // @[Mux.scala 19:72:@31168.4]
  wire [7:0] _T_60947; // @[Mux.scala 19:72:@31175.4]
  wire [15:0] _T_60948; // @[Mux.scala 19:72:@31176.4]
  wire [15:0] _T_60950; // @[Mux.scala 19:72:@31177.4]
  wire [7:0] _T_60957; // @[Mux.scala 19:72:@31184.4]
  wire [7:0] _T_60964; // @[Mux.scala 19:72:@31191.4]
  wire [15:0] _T_60965; // @[Mux.scala 19:72:@31192.4]
  wire [15:0] _T_60967; // @[Mux.scala 19:72:@31193.4]
  wire [7:0] _T_60974; // @[Mux.scala 19:72:@31200.4]
  wire [7:0] _T_60981; // @[Mux.scala 19:72:@31207.4]
  wire [15:0] _T_60982; // @[Mux.scala 19:72:@31208.4]
  wire [15:0] _T_60984; // @[Mux.scala 19:72:@31209.4]
  wire [7:0] _T_60991; // @[Mux.scala 19:72:@31216.4]
  wire [7:0] _T_60998; // @[Mux.scala 19:72:@31223.4]
  wire [15:0] _T_60999; // @[Mux.scala 19:72:@31224.4]
  wire [15:0] _T_61001; // @[Mux.scala 19:72:@31225.4]
  wire [7:0] _T_61008; // @[Mux.scala 19:72:@31232.4]
  wire [7:0] _T_61015; // @[Mux.scala 19:72:@31239.4]
  wire [15:0] _T_61016; // @[Mux.scala 19:72:@31240.4]
  wire [15:0] _T_61018; // @[Mux.scala 19:72:@31241.4]
  wire [7:0] _T_61025; // @[Mux.scala 19:72:@31248.4]
  wire [7:0] _T_61032; // @[Mux.scala 19:72:@31255.4]
  wire [15:0] _T_61033; // @[Mux.scala 19:72:@31256.4]
  wire [15:0] _T_61035; // @[Mux.scala 19:72:@31257.4]
  wire [15:0] _T_61050; // @[Mux.scala 19:72:@31272.4]
  wire [15:0] _T_61052; // @[Mux.scala 19:72:@31273.4]
  wire [15:0] _T_61067; // @[Mux.scala 19:72:@31288.4]
  wire [15:0] _T_61069; // @[Mux.scala 19:72:@31289.4]
  wire [15:0] _T_61084; // @[Mux.scala 19:72:@31304.4]
  wire [15:0] _T_61086; // @[Mux.scala 19:72:@31305.4]
  wire [15:0] _T_61101; // @[Mux.scala 19:72:@31320.4]
  wire [15:0] _T_61103; // @[Mux.scala 19:72:@31321.4]
  wire [15:0] _T_61118; // @[Mux.scala 19:72:@31336.4]
  wire [15:0] _T_61120; // @[Mux.scala 19:72:@31337.4]
  wire [15:0] _T_61135; // @[Mux.scala 19:72:@31352.4]
  wire [15:0] _T_61137; // @[Mux.scala 19:72:@31353.4]
  wire [15:0] _T_61152; // @[Mux.scala 19:72:@31368.4]
  wire [15:0] _T_61154; // @[Mux.scala 19:72:@31369.4]
  wire [15:0] _T_61169; // @[Mux.scala 19:72:@31384.4]
  wire [15:0] _T_61171; // @[Mux.scala 19:72:@31385.4]
  wire [15:0] _T_61172; // @[Mux.scala 19:72:@31386.4]
  wire [15:0] _T_61173; // @[Mux.scala 19:72:@31387.4]
  wire [15:0] _T_61174; // @[Mux.scala 19:72:@31388.4]
  wire [15:0] _T_61175; // @[Mux.scala 19:72:@31389.4]
  wire [15:0] _T_61176; // @[Mux.scala 19:72:@31390.4]
  wire [15:0] _T_61177; // @[Mux.scala 19:72:@31391.4]
  wire [15:0] _T_61178; // @[Mux.scala 19:72:@31392.4]
  wire [15:0] _T_61179; // @[Mux.scala 19:72:@31393.4]
  wire [15:0] _T_61180; // @[Mux.scala 19:72:@31394.4]
  wire [15:0] _T_61181; // @[Mux.scala 19:72:@31395.4]
  wire [15:0] _T_61182; // @[Mux.scala 19:72:@31396.4]
  wire [15:0] _T_61183; // @[Mux.scala 19:72:@31397.4]
  wire [15:0] _T_61184; // @[Mux.scala 19:72:@31398.4]
  wire [15:0] _T_61185; // @[Mux.scala 19:72:@31399.4]
  wire [15:0] _T_61186; // @[Mux.scala 19:72:@31400.4]
  wire [7:0] _T_61764; // @[Mux.scala 19:72:@31750.4]
  wire [7:0] _T_61771; // @[Mux.scala 19:72:@31757.4]
  wire [15:0] _T_61772; // @[Mux.scala 19:72:@31758.4]
  wire [15:0] _T_61774; // @[Mux.scala 19:72:@31759.4]
  wire [7:0] _T_61781; // @[Mux.scala 19:72:@31766.4]
  wire [7:0] _T_61788; // @[Mux.scala 19:72:@31773.4]
  wire [15:0] _T_61789; // @[Mux.scala 19:72:@31774.4]
  wire [15:0] _T_61791; // @[Mux.scala 19:72:@31775.4]
  wire [7:0] _T_61798; // @[Mux.scala 19:72:@31782.4]
  wire [7:0] _T_61805; // @[Mux.scala 19:72:@31789.4]
  wire [15:0] _T_61806; // @[Mux.scala 19:72:@31790.4]
  wire [15:0] _T_61808; // @[Mux.scala 19:72:@31791.4]
  wire [7:0] _T_61815; // @[Mux.scala 19:72:@31798.4]
  wire [7:0] _T_61822; // @[Mux.scala 19:72:@31805.4]
  wire [15:0] _T_61823; // @[Mux.scala 19:72:@31806.4]
  wire [15:0] _T_61825; // @[Mux.scala 19:72:@31807.4]
  wire [7:0] _T_61832; // @[Mux.scala 19:72:@31814.4]
  wire [7:0] _T_61839; // @[Mux.scala 19:72:@31821.4]
  wire [15:0] _T_61840; // @[Mux.scala 19:72:@31822.4]
  wire [15:0] _T_61842; // @[Mux.scala 19:72:@31823.4]
  wire [7:0] _T_61849; // @[Mux.scala 19:72:@31830.4]
  wire [7:0] _T_61856; // @[Mux.scala 19:72:@31837.4]
  wire [15:0] _T_61857; // @[Mux.scala 19:72:@31838.4]
  wire [15:0] _T_61859; // @[Mux.scala 19:72:@31839.4]
  wire [7:0] _T_61866; // @[Mux.scala 19:72:@31846.4]
  wire [7:0] _T_61873; // @[Mux.scala 19:72:@31853.4]
  wire [15:0] _T_61874; // @[Mux.scala 19:72:@31854.4]
  wire [15:0] _T_61876; // @[Mux.scala 19:72:@31855.4]
  wire [7:0] _T_61883; // @[Mux.scala 19:72:@31862.4]
  wire [7:0] _T_61890; // @[Mux.scala 19:72:@31869.4]
  wire [15:0] _T_61891; // @[Mux.scala 19:72:@31870.4]
  wire [15:0] _T_61893; // @[Mux.scala 19:72:@31871.4]
  wire [15:0] _T_61908; // @[Mux.scala 19:72:@31886.4]
  wire [15:0] _T_61910; // @[Mux.scala 19:72:@31887.4]
  wire [15:0] _T_61925; // @[Mux.scala 19:72:@31902.4]
  wire [15:0] _T_61927; // @[Mux.scala 19:72:@31903.4]
  wire [15:0] _T_61942; // @[Mux.scala 19:72:@31918.4]
  wire [15:0] _T_61944; // @[Mux.scala 19:72:@31919.4]
  wire [15:0] _T_61959; // @[Mux.scala 19:72:@31934.4]
  wire [15:0] _T_61961; // @[Mux.scala 19:72:@31935.4]
  wire [15:0] _T_61976; // @[Mux.scala 19:72:@31950.4]
  wire [15:0] _T_61978; // @[Mux.scala 19:72:@31951.4]
  wire [15:0] _T_61993; // @[Mux.scala 19:72:@31966.4]
  wire [15:0] _T_61995; // @[Mux.scala 19:72:@31967.4]
  wire [15:0] _T_62010; // @[Mux.scala 19:72:@31982.4]
  wire [15:0] _T_62012; // @[Mux.scala 19:72:@31983.4]
  wire [15:0] _T_62027; // @[Mux.scala 19:72:@31998.4]
  wire [15:0] _T_62029; // @[Mux.scala 19:72:@31999.4]
  wire [15:0] _T_62030; // @[Mux.scala 19:72:@32000.4]
  wire [15:0] _T_62031; // @[Mux.scala 19:72:@32001.4]
  wire [15:0] _T_62032; // @[Mux.scala 19:72:@32002.4]
  wire [15:0] _T_62033; // @[Mux.scala 19:72:@32003.4]
  wire [15:0] _T_62034; // @[Mux.scala 19:72:@32004.4]
  wire [15:0] _T_62035; // @[Mux.scala 19:72:@32005.4]
  wire [15:0] _T_62036; // @[Mux.scala 19:72:@32006.4]
  wire [15:0] _T_62037; // @[Mux.scala 19:72:@32007.4]
  wire [15:0] _T_62038; // @[Mux.scala 19:72:@32008.4]
  wire [15:0] _T_62039; // @[Mux.scala 19:72:@32009.4]
  wire [15:0] _T_62040; // @[Mux.scala 19:72:@32010.4]
  wire [15:0] _T_62041; // @[Mux.scala 19:72:@32011.4]
  wire [15:0] _T_62042; // @[Mux.scala 19:72:@32012.4]
  wire [15:0] _T_62043; // @[Mux.scala 19:72:@32013.4]
  wire [15:0] _T_62044; // @[Mux.scala 19:72:@32014.4]
  wire [7:0] _T_62622; // @[Mux.scala 19:72:@32364.4]
  wire [7:0] _T_62629; // @[Mux.scala 19:72:@32371.4]
  wire [15:0] _T_62630; // @[Mux.scala 19:72:@32372.4]
  wire [15:0] _T_62632; // @[Mux.scala 19:72:@32373.4]
  wire [7:0] _T_62639; // @[Mux.scala 19:72:@32380.4]
  wire [7:0] _T_62646; // @[Mux.scala 19:72:@32387.4]
  wire [15:0] _T_62647; // @[Mux.scala 19:72:@32388.4]
  wire [15:0] _T_62649; // @[Mux.scala 19:72:@32389.4]
  wire [7:0] _T_62656; // @[Mux.scala 19:72:@32396.4]
  wire [7:0] _T_62663; // @[Mux.scala 19:72:@32403.4]
  wire [15:0] _T_62664; // @[Mux.scala 19:72:@32404.4]
  wire [15:0] _T_62666; // @[Mux.scala 19:72:@32405.4]
  wire [7:0] _T_62673; // @[Mux.scala 19:72:@32412.4]
  wire [7:0] _T_62680; // @[Mux.scala 19:72:@32419.4]
  wire [15:0] _T_62681; // @[Mux.scala 19:72:@32420.4]
  wire [15:0] _T_62683; // @[Mux.scala 19:72:@32421.4]
  wire [7:0] _T_62690; // @[Mux.scala 19:72:@32428.4]
  wire [7:0] _T_62697; // @[Mux.scala 19:72:@32435.4]
  wire [15:0] _T_62698; // @[Mux.scala 19:72:@32436.4]
  wire [15:0] _T_62700; // @[Mux.scala 19:72:@32437.4]
  wire [7:0] _T_62707; // @[Mux.scala 19:72:@32444.4]
  wire [7:0] _T_62714; // @[Mux.scala 19:72:@32451.4]
  wire [15:0] _T_62715; // @[Mux.scala 19:72:@32452.4]
  wire [15:0] _T_62717; // @[Mux.scala 19:72:@32453.4]
  wire [7:0] _T_62724; // @[Mux.scala 19:72:@32460.4]
  wire [7:0] _T_62731; // @[Mux.scala 19:72:@32467.4]
  wire [15:0] _T_62732; // @[Mux.scala 19:72:@32468.4]
  wire [15:0] _T_62734; // @[Mux.scala 19:72:@32469.4]
  wire [7:0] _T_62741; // @[Mux.scala 19:72:@32476.4]
  wire [7:0] _T_62748; // @[Mux.scala 19:72:@32483.4]
  wire [15:0] _T_62749; // @[Mux.scala 19:72:@32484.4]
  wire [15:0] _T_62751; // @[Mux.scala 19:72:@32485.4]
  wire [15:0] _T_62766; // @[Mux.scala 19:72:@32500.4]
  wire [15:0] _T_62768; // @[Mux.scala 19:72:@32501.4]
  wire [15:0] _T_62783; // @[Mux.scala 19:72:@32516.4]
  wire [15:0] _T_62785; // @[Mux.scala 19:72:@32517.4]
  wire [15:0] _T_62800; // @[Mux.scala 19:72:@32532.4]
  wire [15:0] _T_62802; // @[Mux.scala 19:72:@32533.4]
  wire [15:0] _T_62817; // @[Mux.scala 19:72:@32548.4]
  wire [15:0] _T_62819; // @[Mux.scala 19:72:@32549.4]
  wire [15:0] _T_62834; // @[Mux.scala 19:72:@32564.4]
  wire [15:0] _T_62836; // @[Mux.scala 19:72:@32565.4]
  wire [15:0] _T_62851; // @[Mux.scala 19:72:@32580.4]
  wire [15:0] _T_62853; // @[Mux.scala 19:72:@32581.4]
  wire [15:0] _T_62868; // @[Mux.scala 19:72:@32596.4]
  wire [15:0] _T_62870; // @[Mux.scala 19:72:@32597.4]
  wire [15:0] _T_62885; // @[Mux.scala 19:72:@32612.4]
  wire [15:0] _T_62887; // @[Mux.scala 19:72:@32613.4]
  wire [15:0] _T_62888; // @[Mux.scala 19:72:@32614.4]
  wire [15:0] _T_62889; // @[Mux.scala 19:72:@32615.4]
  wire [15:0] _T_62890; // @[Mux.scala 19:72:@32616.4]
  wire [15:0] _T_62891; // @[Mux.scala 19:72:@32617.4]
  wire [15:0] _T_62892; // @[Mux.scala 19:72:@32618.4]
  wire [15:0] _T_62893; // @[Mux.scala 19:72:@32619.4]
  wire [15:0] _T_62894; // @[Mux.scala 19:72:@32620.4]
  wire [15:0] _T_62895; // @[Mux.scala 19:72:@32621.4]
  wire [15:0] _T_62896; // @[Mux.scala 19:72:@32622.4]
  wire [15:0] _T_62897; // @[Mux.scala 19:72:@32623.4]
  wire [15:0] _T_62898; // @[Mux.scala 19:72:@32624.4]
  wire [15:0] _T_62899; // @[Mux.scala 19:72:@32625.4]
  wire [15:0] _T_62900; // @[Mux.scala 19:72:@32626.4]
  wire [15:0] _T_62901; // @[Mux.scala 19:72:@32627.4]
  wire [15:0] _T_62902; // @[Mux.scala 19:72:@32628.4]
  wire [7:0] _T_63480; // @[Mux.scala 19:72:@32978.4]
  wire [7:0] _T_63487; // @[Mux.scala 19:72:@32985.4]
  wire [15:0] _T_63488; // @[Mux.scala 19:72:@32986.4]
  wire [15:0] _T_63490; // @[Mux.scala 19:72:@32987.4]
  wire [7:0] _T_63497; // @[Mux.scala 19:72:@32994.4]
  wire [7:0] _T_63504; // @[Mux.scala 19:72:@33001.4]
  wire [15:0] _T_63505; // @[Mux.scala 19:72:@33002.4]
  wire [15:0] _T_63507; // @[Mux.scala 19:72:@33003.4]
  wire [7:0] _T_63514; // @[Mux.scala 19:72:@33010.4]
  wire [7:0] _T_63521; // @[Mux.scala 19:72:@33017.4]
  wire [15:0] _T_63522; // @[Mux.scala 19:72:@33018.4]
  wire [15:0] _T_63524; // @[Mux.scala 19:72:@33019.4]
  wire [7:0] _T_63531; // @[Mux.scala 19:72:@33026.4]
  wire [7:0] _T_63538; // @[Mux.scala 19:72:@33033.4]
  wire [15:0] _T_63539; // @[Mux.scala 19:72:@33034.4]
  wire [15:0] _T_63541; // @[Mux.scala 19:72:@33035.4]
  wire [7:0] _T_63548; // @[Mux.scala 19:72:@33042.4]
  wire [7:0] _T_63555; // @[Mux.scala 19:72:@33049.4]
  wire [15:0] _T_63556; // @[Mux.scala 19:72:@33050.4]
  wire [15:0] _T_63558; // @[Mux.scala 19:72:@33051.4]
  wire [7:0] _T_63565; // @[Mux.scala 19:72:@33058.4]
  wire [7:0] _T_63572; // @[Mux.scala 19:72:@33065.4]
  wire [15:0] _T_63573; // @[Mux.scala 19:72:@33066.4]
  wire [15:0] _T_63575; // @[Mux.scala 19:72:@33067.4]
  wire [7:0] _T_63582; // @[Mux.scala 19:72:@33074.4]
  wire [7:0] _T_63589; // @[Mux.scala 19:72:@33081.4]
  wire [15:0] _T_63590; // @[Mux.scala 19:72:@33082.4]
  wire [15:0] _T_63592; // @[Mux.scala 19:72:@33083.4]
  wire [7:0] _T_63599; // @[Mux.scala 19:72:@33090.4]
  wire [7:0] _T_63606; // @[Mux.scala 19:72:@33097.4]
  wire [15:0] _T_63607; // @[Mux.scala 19:72:@33098.4]
  wire [15:0] _T_63609; // @[Mux.scala 19:72:@33099.4]
  wire [15:0] _T_63624; // @[Mux.scala 19:72:@33114.4]
  wire [15:0] _T_63626; // @[Mux.scala 19:72:@33115.4]
  wire [15:0] _T_63641; // @[Mux.scala 19:72:@33130.4]
  wire [15:0] _T_63643; // @[Mux.scala 19:72:@33131.4]
  wire [15:0] _T_63658; // @[Mux.scala 19:72:@33146.4]
  wire [15:0] _T_63660; // @[Mux.scala 19:72:@33147.4]
  wire [15:0] _T_63675; // @[Mux.scala 19:72:@33162.4]
  wire [15:0] _T_63677; // @[Mux.scala 19:72:@33163.4]
  wire [15:0] _T_63692; // @[Mux.scala 19:72:@33178.4]
  wire [15:0] _T_63694; // @[Mux.scala 19:72:@33179.4]
  wire [15:0] _T_63709; // @[Mux.scala 19:72:@33194.4]
  wire [15:0] _T_63711; // @[Mux.scala 19:72:@33195.4]
  wire [15:0] _T_63726; // @[Mux.scala 19:72:@33210.4]
  wire [15:0] _T_63728; // @[Mux.scala 19:72:@33211.4]
  wire [15:0] _T_63743; // @[Mux.scala 19:72:@33226.4]
  wire [15:0] _T_63745; // @[Mux.scala 19:72:@33227.4]
  wire [15:0] _T_63746; // @[Mux.scala 19:72:@33228.4]
  wire [15:0] _T_63747; // @[Mux.scala 19:72:@33229.4]
  wire [15:0] _T_63748; // @[Mux.scala 19:72:@33230.4]
  wire [15:0] _T_63749; // @[Mux.scala 19:72:@33231.4]
  wire [15:0] _T_63750; // @[Mux.scala 19:72:@33232.4]
  wire [15:0] _T_63751; // @[Mux.scala 19:72:@33233.4]
  wire [15:0] _T_63752; // @[Mux.scala 19:72:@33234.4]
  wire [15:0] _T_63753; // @[Mux.scala 19:72:@33235.4]
  wire [15:0] _T_63754; // @[Mux.scala 19:72:@33236.4]
  wire [15:0] _T_63755; // @[Mux.scala 19:72:@33237.4]
  wire [15:0] _T_63756; // @[Mux.scala 19:72:@33238.4]
  wire [15:0] _T_63757; // @[Mux.scala 19:72:@33239.4]
  wire [15:0] _T_63758; // @[Mux.scala 19:72:@33240.4]
  wire [15:0] _T_63759; // @[Mux.scala 19:72:@33241.4]
  wire [15:0] _T_63760; // @[Mux.scala 19:72:@33242.4]
  wire [7:0] _T_64338; // @[Mux.scala 19:72:@33592.4]
  wire [7:0] _T_64345; // @[Mux.scala 19:72:@33599.4]
  wire [15:0] _T_64346; // @[Mux.scala 19:72:@33600.4]
  wire [15:0] _T_64348; // @[Mux.scala 19:72:@33601.4]
  wire [7:0] _T_64355; // @[Mux.scala 19:72:@33608.4]
  wire [7:0] _T_64362; // @[Mux.scala 19:72:@33615.4]
  wire [15:0] _T_64363; // @[Mux.scala 19:72:@33616.4]
  wire [15:0] _T_64365; // @[Mux.scala 19:72:@33617.4]
  wire [7:0] _T_64372; // @[Mux.scala 19:72:@33624.4]
  wire [7:0] _T_64379; // @[Mux.scala 19:72:@33631.4]
  wire [15:0] _T_64380; // @[Mux.scala 19:72:@33632.4]
  wire [15:0] _T_64382; // @[Mux.scala 19:72:@33633.4]
  wire [7:0] _T_64389; // @[Mux.scala 19:72:@33640.4]
  wire [7:0] _T_64396; // @[Mux.scala 19:72:@33647.4]
  wire [15:0] _T_64397; // @[Mux.scala 19:72:@33648.4]
  wire [15:0] _T_64399; // @[Mux.scala 19:72:@33649.4]
  wire [7:0] _T_64406; // @[Mux.scala 19:72:@33656.4]
  wire [7:0] _T_64413; // @[Mux.scala 19:72:@33663.4]
  wire [15:0] _T_64414; // @[Mux.scala 19:72:@33664.4]
  wire [15:0] _T_64416; // @[Mux.scala 19:72:@33665.4]
  wire [7:0] _T_64423; // @[Mux.scala 19:72:@33672.4]
  wire [7:0] _T_64430; // @[Mux.scala 19:72:@33679.4]
  wire [15:0] _T_64431; // @[Mux.scala 19:72:@33680.4]
  wire [15:0] _T_64433; // @[Mux.scala 19:72:@33681.4]
  wire [7:0] _T_64440; // @[Mux.scala 19:72:@33688.4]
  wire [7:0] _T_64447; // @[Mux.scala 19:72:@33695.4]
  wire [15:0] _T_64448; // @[Mux.scala 19:72:@33696.4]
  wire [15:0] _T_64450; // @[Mux.scala 19:72:@33697.4]
  wire [7:0] _T_64457; // @[Mux.scala 19:72:@33704.4]
  wire [7:0] _T_64464; // @[Mux.scala 19:72:@33711.4]
  wire [15:0] _T_64465; // @[Mux.scala 19:72:@33712.4]
  wire [15:0] _T_64467; // @[Mux.scala 19:72:@33713.4]
  wire [15:0] _T_64482; // @[Mux.scala 19:72:@33728.4]
  wire [15:0] _T_64484; // @[Mux.scala 19:72:@33729.4]
  wire [15:0] _T_64499; // @[Mux.scala 19:72:@33744.4]
  wire [15:0] _T_64501; // @[Mux.scala 19:72:@33745.4]
  wire [15:0] _T_64516; // @[Mux.scala 19:72:@33760.4]
  wire [15:0] _T_64518; // @[Mux.scala 19:72:@33761.4]
  wire [15:0] _T_64533; // @[Mux.scala 19:72:@33776.4]
  wire [15:0] _T_64535; // @[Mux.scala 19:72:@33777.4]
  wire [15:0] _T_64550; // @[Mux.scala 19:72:@33792.4]
  wire [15:0] _T_64552; // @[Mux.scala 19:72:@33793.4]
  wire [15:0] _T_64567; // @[Mux.scala 19:72:@33808.4]
  wire [15:0] _T_64569; // @[Mux.scala 19:72:@33809.4]
  wire [15:0] _T_64584; // @[Mux.scala 19:72:@33824.4]
  wire [15:0] _T_64586; // @[Mux.scala 19:72:@33825.4]
  wire [15:0] _T_64601; // @[Mux.scala 19:72:@33840.4]
  wire [15:0] _T_64603; // @[Mux.scala 19:72:@33841.4]
  wire [15:0] _T_64604; // @[Mux.scala 19:72:@33842.4]
  wire [15:0] _T_64605; // @[Mux.scala 19:72:@33843.4]
  wire [15:0] _T_64606; // @[Mux.scala 19:72:@33844.4]
  wire [15:0] _T_64607; // @[Mux.scala 19:72:@33845.4]
  wire [15:0] _T_64608; // @[Mux.scala 19:72:@33846.4]
  wire [15:0] _T_64609; // @[Mux.scala 19:72:@33847.4]
  wire [15:0] _T_64610; // @[Mux.scala 19:72:@33848.4]
  wire [15:0] _T_64611; // @[Mux.scala 19:72:@33849.4]
  wire [15:0] _T_64612; // @[Mux.scala 19:72:@33850.4]
  wire [15:0] _T_64613; // @[Mux.scala 19:72:@33851.4]
  wire [15:0] _T_64614; // @[Mux.scala 19:72:@33852.4]
  wire [15:0] _T_64615; // @[Mux.scala 19:72:@33853.4]
  wire [15:0] _T_64616; // @[Mux.scala 19:72:@33854.4]
  wire [15:0] _T_64617; // @[Mux.scala 19:72:@33855.4]
  wire [15:0] _T_64618; // @[Mux.scala 19:72:@33856.4]
  wire [7:0] _T_65196; // @[Mux.scala 19:72:@34206.4]
  wire [7:0] _T_65203; // @[Mux.scala 19:72:@34213.4]
  wire [15:0] _T_65204; // @[Mux.scala 19:72:@34214.4]
  wire [15:0] _T_65206; // @[Mux.scala 19:72:@34215.4]
  wire [7:0] _T_65213; // @[Mux.scala 19:72:@34222.4]
  wire [7:0] _T_65220; // @[Mux.scala 19:72:@34229.4]
  wire [15:0] _T_65221; // @[Mux.scala 19:72:@34230.4]
  wire [15:0] _T_65223; // @[Mux.scala 19:72:@34231.4]
  wire [7:0] _T_65230; // @[Mux.scala 19:72:@34238.4]
  wire [7:0] _T_65237; // @[Mux.scala 19:72:@34245.4]
  wire [15:0] _T_65238; // @[Mux.scala 19:72:@34246.4]
  wire [15:0] _T_65240; // @[Mux.scala 19:72:@34247.4]
  wire [7:0] _T_65247; // @[Mux.scala 19:72:@34254.4]
  wire [7:0] _T_65254; // @[Mux.scala 19:72:@34261.4]
  wire [15:0] _T_65255; // @[Mux.scala 19:72:@34262.4]
  wire [15:0] _T_65257; // @[Mux.scala 19:72:@34263.4]
  wire [7:0] _T_65264; // @[Mux.scala 19:72:@34270.4]
  wire [7:0] _T_65271; // @[Mux.scala 19:72:@34277.4]
  wire [15:0] _T_65272; // @[Mux.scala 19:72:@34278.4]
  wire [15:0] _T_65274; // @[Mux.scala 19:72:@34279.4]
  wire [7:0] _T_65281; // @[Mux.scala 19:72:@34286.4]
  wire [7:0] _T_65288; // @[Mux.scala 19:72:@34293.4]
  wire [15:0] _T_65289; // @[Mux.scala 19:72:@34294.4]
  wire [15:0] _T_65291; // @[Mux.scala 19:72:@34295.4]
  wire [7:0] _T_65298; // @[Mux.scala 19:72:@34302.4]
  wire [7:0] _T_65305; // @[Mux.scala 19:72:@34309.4]
  wire [15:0] _T_65306; // @[Mux.scala 19:72:@34310.4]
  wire [15:0] _T_65308; // @[Mux.scala 19:72:@34311.4]
  wire [7:0] _T_65315; // @[Mux.scala 19:72:@34318.4]
  wire [7:0] _T_65322; // @[Mux.scala 19:72:@34325.4]
  wire [15:0] _T_65323; // @[Mux.scala 19:72:@34326.4]
  wire [15:0] _T_65325; // @[Mux.scala 19:72:@34327.4]
  wire [15:0] _T_65340; // @[Mux.scala 19:72:@34342.4]
  wire [15:0] _T_65342; // @[Mux.scala 19:72:@34343.4]
  wire [15:0] _T_65357; // @[Mux.scala 19:72:@34358.4]
  wire [15:0] _T_65359; // @[Mux.scala 19:72:@34359.4]
  wire [15:0] _T_65374; // @[Mux.scala 19:72:@34374.4]
  wire [15:0] _T_65376; // @[Mux.scala 19:72:@34375.4]
  wire [15:0] _T_65391; // @[Mux.scala 19:72:@34390.4]
  wire [15:0] _T_65393; // @[Mux.scala 19:72:@34391.4]
  wire [15:0] _T_65408; // @[Mux.scala 19:72:@34406.4]
  wire [15:0] _T_65410; // @[Mux.scala 19:72:@34407.4]
  wire [15:0] _T_65425; // @[Mux.scala 19:72:@34422.4]
  wire [15:0] _T_65427; // @[Mux.scala 19:72:@34423.4]
  wire [15:0] _T_65442; // @[Mux.scala 19:72:@34438.4]
  wire [15:0] _T_65444; // @[Mux.scala 19:72:@34439.4]
  wire [15:0] _T_65459; // @[Mux.scala 19:72:@34454.4]
  wire [15:0] _T_65461; // @[Mux.scala 19:72:@34455.4]
  wire [15:0] _T_65462; // @[Mux.scala 19:72:@34456.4]
  wire [15:0] _T_65463; // @[Mux.scala 19:72:@34457.4]
  wire [15:0] _T_65464; // @[Mux.scala 19:72:@34458.4]
  wire [15:0] _T_65465; // @[Mux.scala 19:72:@34459.4]
  wire [15:0] _T_65466; // @[Mux.scala 19:72:@34460.4]
  wire [15:0] _T_65467; // @[Mux.scala 19:72:@34461.4]
  wire [15:0] _T_65468; // @[Mux.scala 19:72:@34462.4]
  wire [15:0] _T_65469; // @[Mux.scala 19:72:@34463.4]
  wire [15:0] _T_65470; // @[Mux.scala 19:72:@34464.4]
  wire [15:0] _T_65471; // @[Mux.scala 19:72:@34465.4]
  wire [15:0] _T_65472; // @[Mux.scala 19:72:@34466.4]
  wire [15:0] _T_65473; // @[Mux.scala 19:72:@34467.4]
  wire [15:0] _T_65474; // @[Mux.scala 19:72:@34468.4]
  wire [15:0] _T_65475; // @[Mux.scala 19:72:@34469.4]
  wire [15:0] _T_65476; // @[Mux.scala 19:72:@34470.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_419;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_420;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_421;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_422;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_423;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_424;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_425;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_426;
  reg  storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_427;
  reg  storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_428;
  reg  storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_429;
  reg  storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_430;
  reg  storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_431;
  reg  storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_432;
  reg  storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_433;
  reg  storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_434;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_435;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_436;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_437;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_438;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_439;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_440;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_441;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_442;
  reg  storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_443;
  reg  storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_444;
  reg  storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_445;
  reg  storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_446;
  reg  storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_447;
  reg  storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_448;
  reg  storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_449;
  reg  storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_450;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_451;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_452;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_453;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_454;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_455;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_456;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_457;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_458;
  reg  storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_459;
  reg  storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_460;
  reg  storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_461;
  reg  storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_462;
  reg  storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_463;
  reg  storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_464;
  reg  storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_465;
  reg  storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_466;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_467;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_468;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_469;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_470;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_471;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_472;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_473;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_474;
  reg  storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_475;
  reg  storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_476;
  reg  storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_477;
  reg  storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_478;
  reg  storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_479;
  reg  storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_480;
  reg  storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_481;
  reg  storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_482;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_483;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_484;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_485;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_486;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_487;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_488;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_489;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_490;
  reg  storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_491;
  reg  storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_492;
  reg  storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_493;
  reg  storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_494;
  reg  storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_495;
  reg  storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_496;
  reg  storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_497;
  reg  storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_498;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_499;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_500;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_501;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_502;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_503;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_504;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_505;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_506;
  reg  storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_507;
  reg  storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_508;
  reg  storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_509;
  reg  storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_510;
  reg  storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_511;
  reg  storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_512;
  reg  storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_513;
  reg  storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_514;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_515;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_516;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_517;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_518;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_519;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_520;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_521;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_522;
  reg  storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_523;
  reg  storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_524;
  reg  storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_525;
  reg  storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_526;
  reg  storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_527;
  reg  storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_528;
  reg  storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_529;
  reg  storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_530;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_531;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_532;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_533;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_534;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_535;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_536;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_537;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_538;
  reg  storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_539;
  reg  storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_540;
  reg  storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_541;
  reg  storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_542;
  reg  storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_543;
  reg  storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_544;
  reg  storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_545;
  reg  storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_546;
  reg  storeAddrNotKnownFlagsPReg_8_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_547;
  reg  storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_548;
  reg  storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_549;
  reg  storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_550;
  reg  storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_551;
  reg  storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_552;
  reg  storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_553;
  reg  storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_554;
  reg  storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_555;
  reg  storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_556;
  reg  storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_557;
  reg  storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_558;
  reg  storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_559;
  reg  storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_560;
  reg  storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_561;
  reg  storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_562;
  reg  storeAddrNotKnownFlagsPReg_9_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_563;
  reg  storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_564;
  reg  storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_565;
  reg  storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_566;
  reg  storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_567;
  reg  storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_568;
  reg  storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_569;
  reg  storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_570;
  reg  storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_571;
  reg  storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_572;
  reg  storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_573;
  reg  storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_574;
  reg  storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_575;
  reg  storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_576;
  reg  storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_577;
  reg  storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_578;
  reg  storeAddrNotKnownFlagsPReg_10_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_579;
  reg  storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_580;
  reg  storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_581;
  reg  storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_582;
  reg  storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_583;
  reg  storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_584;
  reg  storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_585;
  reg  storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_586;
  reg  storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_587;
  reg  storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_588;
  reg  storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_589;
  reg  storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_590;
  reg  storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_591;
  reg  storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_592;
  reg  storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_593;
  reg  storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_594;
  reg  storeAddrNotKnownFlagsPReg_11_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_595;
  reg  storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_596;
  reg  storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_597;
  reg  storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_598;
  reg  storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_599;
  reg  storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_600;
  reg  storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_601;
  reg  storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_602;
  reg  storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_603;
  reg  storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_604;
  reg  storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_605;
  reg  storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_606;
  reg  storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_607;
  reg  storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_608;
  reg  storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_609;
  reg  storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_610;
  reg  storeAddrNotKnownFlagsPReg_12_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_611;
  reg  storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_612;
  reg  storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_613;
  reg  storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_614;
  reg  storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_615;
  reg  storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_616;
  reg  storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_617;
  reg  storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_618;
  reg  storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_619;
  reg  storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_620;
  reg  storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_621;
  reg  storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_622;
  reg  storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_623;
  reg  storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_624;
  reg  storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_625;
  reg  storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_626;
  reg  storeAddrNotKnownFlagsPReg_13_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_627;
  reg  storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_628;
  reg  storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_629;
  reg  storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_630;
  reg  storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_631;
  reg  storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_632;
  reg  storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_633;
  reg  storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_634;
  reg  storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_635;
  reg  storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_636;
  reg  storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_637;
  reg  storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_638;
  reg  storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_639;
  reg  storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_640;
  reg  storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_641;
  reg  storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_642;
  reg  storeAddrNotKnownFlagsPReg_14_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_643;
  reg  storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_644;
  reg  storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_645;
  reg  storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_646;
  reg  storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_647;
  reg  storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_648;
  reg  storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_649;
  reg  storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_650;
  reg  storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_651;
  reg  storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_652;
  reg  storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_653;
  reg  storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_654;
  reg  storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_655;
  reg  storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_656;
  reg  storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_657;
  reg  storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_658;
  reg  storeAddrNotKnownFlagsPReg_15_0; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_659;
  reg  storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_660;
  reg  storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_661;
  reg  storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_662;
  reg  storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_663;
  reg  storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_664;
  reg  storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_665;
  reg  storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_666;
  reg  storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_667;
  reg  storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_668;
  reg  storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_669;
  reg  storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_670;
  reg  storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_671;
  reg  storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_672;
  reg  storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_673;
  reg  storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 167:43:@34763.4]
  reg [31:0] _RAND_674;
  reg  shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_675;
  reg  shiftedStoreDataKnownPReg_1; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_676;
  reg  shiftedStoreDataKnownPReg_2; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_677;
  reg  shiftedStoreDataKnownPReg_3; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_678;
  reg  shiftedStoreDataKnownPReg_4; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_679;
  reg  shiftedStoreDataKnownPReg_5; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_680;
  reg  shiftedStoreDataKnownPReg_6; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_681;
  reg  shiftedStoreDataKnownPReg_7; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_682;
  reg  shiftedStoreDataKnownPReg_8; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_683;
  reg  shiftedStoreDataKnownPReg_9; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_684;
  reg  shiftedStoreDataKnownPReg_10; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_685;
  reg  shiftedStoreDataKnownPReg_11; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_686;
  reg  shiftedStoreDataKnownPReg_12; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_687;
  reg  shiftedStoreDataKnownPReg_13; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_688;
  reg  shiftedStoreDataKnownPReg_14; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_689;
  reg  shiftedStoreDataKnownPReg_15; // @[LoadQueue.scala 168:42:@35020.4]
  reg [31:0] _RAND_690;
  reg [31:0] shiftedStoreDataQPreg_0; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_691;
  reg [31:0] shiftedStoreDataQPreg_1; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_692;
  reg [31:0] shiftedStoreDataQPreg_2; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_693;
  reg [31:0] shiftedStoreDataQPreg_3; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_694;
  reg [31:0] shiftedStoreDataQPreg_4; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_695;
  reg [31:0] shiftedStoreDataQPreg_5; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_696;
  reg [31:0] shiftedStoreDataQPreg_6; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_697;
  reg [31:0] shiftedStoreDataQPreg_7; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_698;
  reg [31:0] shiftedStoreDataQPreg_8; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_699;
  reg [31:0] shiftedStoreDataQPreg_9; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_700;
  reg [31:0] shiftedStoreDataQPreg_10; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_701;
  reg [31:0] shiftedStoreDataQPreg_11; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_702;
  reg [31:0] shiftedStoreDataQPreg_12; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_703;
  reg [31:0] shiftedStoreDataQPreg_13; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_704;
  reg [31:0] shiftedStoreDataQPreg_14; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_705;
  reg [31:0] shiftedStoreDataQPreg_15; // @[LoadQueue.scala 169:38:@35037.4]
  reg [31:0] _RAND_706;
  reg  addrKnownPReg_0; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_707;
  reg  addrKnownPReg_1; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_708;
  reg  addrKnownPReg_2; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_709;
  reg  addrKnownPReg_3; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_710;
  reg  addrKnownPReg_4; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_711;
  reg  addrKnownPReg_5; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_712;
  reg  addrKnownPReg_6; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_713;
  reg  addrKnownPReg_7; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_714;
  reg  addrKnownPReg_8; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_715;
  reg  addrKnownPReg_9; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_716;
  reg  addrKnownPReg_10; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_717;
  reg  addrKnownPReg_11; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_718;
  reg  addrKnownPReg_12; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_719;
  reg  addrKnownPReg_13; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_720;
  reg  addrKnownPReg_14; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_721;
  reg  addrKnownPReg_15; // @[LoadQueue.scala 170:30:@35054.4]
  reg [31:0] _RAND_722;
  reg  dataKnownPReg_0; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_723;
  reg  dataKnownPReg_1; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_724;
  reg  dataKnownPReg_2; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_725;
  reg  dataKnownPReg_3; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_726;
  reg  dataKnownPReg_4; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_727;
  reg  dataKnownPReg_5; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_728;
  reg  dataKnownPReg_6; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_729;
  reg  dataKnownPReg_7; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_730;
  reg  dataKnownPReg_8; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_731;
  reg  dataKnownPReg_9; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_732;
  reg  dataKnownPReg_10; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_733;
  reg  dataKnownPReg_11; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_734;
  reg  dataKnownPReg_12; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_735;
  reg  dataKnownPReg_13; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_736;
  reg  dataKnownPReg_14; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_737;
  reg  dataKnownPReg_15; // @[LoadQueue.scala 171:30:@35071.4]
  reg [31:0] _RAND_738;
  wire [1:0] _T_88268; // @[LoadQueue.scala 191:60:@35143.4]
  wire [1:0] _T_88269; // @[LoadQueue.scala 191:60:@35144.4]
  wire [2:0] _T_88270; // @[LoadQueue.scala 191:60:@35145.4]
  wire [2:0] _T_88271; // @[LoadQueue.scala 191:60:@35146.4]
  wire [2:0] _T_88272; // @[LoadQueue.scala 191:60:@35147.4]
  wire [2:0] _T_88273; // @[LoadQueue.scala 191:60:@35148.4]
  wire [3:0] _T_88274; // @[LoadQueue.scala 191:60:@35149.4]
  wire [3:0] _T_88275; // @[LoadQueue.scala 191:60:@35150.4]
  wire [3:0] _T_88276; // @[LoadQueue.scala 191:60:@35151.4]
  wire [3:0] _T_88277; // @[LoadQueue.scala 191:60:@35152.4]
  wire [3:0] _T_88278; // @[LoadQueue.scala 191:60:@35153.4]
  wire [3:0] _T_88279; // @[LoadQueue.scala 191:60:@35154.4]
  wire [3:0] _T_88280; // @[LoadQueue.scala 191:60:@35155.4]
  wire [3:0] _T_88281; // @[LoadQueue.scala 191:60:@35156.4]
  wire  _T_88284; // @[LoadQueue.scala 192:43:@35158.4]
  wire  _T_88285; // @[LoadQueue.scala 192:43:@35159.4]
  wire  _T_88286; // @[LoadQueue.scala 192:43:@35160.4]
  wire  _T_88287; // @[LoadQueue.scala 192:43:@35161.4]
  wire  _T_88288; // @[LoadQueue.scala 192:43:@35162.4]
  wire  _T_88289; // @[LoadQueue.scala 192:43:@35163.4]
  wire  _T_88290; // @[LoadQueue.scala 192:43:@35164.4]
  wire  _T_88291; // @[LoadQueue.scala 192:43:@35165.4]
  wire  _T_88292; // @[LoadQueue.scala 192:43:@35166.4]
  wire  _T_88293; // @[LoadQueue.scala 192:43:@35167.4]
  wire  _T_88294; // @[LoadQueue.scala 192:43:@35168.4]
  wire  _T_88295; // @[LoadQueue.scala 192:43:@35169.4]
  wire  _T_88296; // @[LoadQueue.scala 192:43:@35170.4]
  wire  _T_88297; // @[LoadQueue.scala 192:43:@35171.4]
  wire  _T_88298; // @[LoadQueue.scala 192:43:@35172.4]
  wire  _GEN_864; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_865; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_866; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_867; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_868; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_869; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_870; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_871; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_872; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_873; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_874; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_875; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_876; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_877; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_878; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_879; // @[LoadQueue.scala 193:43:@35174.6]
  wire  _GEN_881; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_882; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_883; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_884; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_885; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_886; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_887; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_888; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_889; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_890; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_891; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_892; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_893; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_894; // @[LoadQueue.scala 194:31:@35175.6]
  wire  _GEN_895; // @[LoadQueue.scala 194:31:@35175.6]
  wire [31:0] _GEN_897; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_898; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_899; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_900; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_901; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_902; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_903; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_904; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_905; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_906; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_907; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_908; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_909; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_910; // @[LoadQueue.scala 195:31:@35176.6]
  wire [31:0] _GEN_911; // @[LoadQueue.scala 195:31:@35176.6]
  wire  lastConflict_0_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_1; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_2; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_3; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_4; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_5; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_6; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_7; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_8; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_9; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_10; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_11; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_12; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_13; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_14; // @[LoadQueue.scala 192:53:@35173.4]
  wire  lastConflict_0_15; // @[LoadQueue.scala 192:53:@35173.4]
  wire  canBypass_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire [31:0] bypassVal_0; // @[LoadQueue.scala 192:53:@35173.4]
  wire [1:0] _T_88404; // @[LoadQueue.scala 191:60:@35230.4]
  wire [1:0] _T_88405; // @[LoadQueue.scala 191:60:@35231.4]
  wire [2:0] _T_88406; // @[LoadQueue.scala 191:60:@35232.4]
  wire [2:0] _T_88407; // @[LoadQueue.scala 191:60:@35233.4]
  wire [2:0] _T_88408; // @[LoadQueue.scala 191:60:@35234.4]
  wire [2:0] _T_88409; // @[LoadQueue.scala 191:60:@35235.4]
  wire [3:0] _T_88410; // @[LoadQueue.scala 191:60:@35236.4]
  wire [3:0] _T_88411; // @[LoadQueue.scala 191:60:@35237.4]
  wire [3:0] _T_88412; // @[LoadQueue.scala 191:60:@35238.4]
  wire [3:0] _T_88413; // @[LoadQueue.scala 191:60:@35239.4]
  wire [3:0] _T_88414; // @[LoadQueue.scala 191:60:@35240.4]
  wire [3:0] _T_88415; // @[LoadQueue.scala 191:60:@35241.4]
  wire [3:0] _T_88416; // @[LoadQueue.scala 191:60:@35242.4]
  wire [3:0] _T_88417; // @[LoadQueue.scala 191:60:@35243.4]
  wire  _T_88420; // @[LoadQueue.scala 192:43:@35245.4]
  wire  _T_88421; // @[LoadQueue.scala 192:43:@35246.4]
  wire  _T_88422; // @[LoadQueue.scala 192:43:@35247.4]
  wire  _T_88423; // @[LoadQueue.scala 192:43:@35248.4]
  wire  _T_88424; // @[LoadQueue.scala 192:43:@35249.4]
  wire  _T_88425; // @[LoadQueue.scala 192:43:@35250.4]
  wire  _T_88426; // @[LoadQueue.scala 192:43:@35251.4]
  wire  _T_88427; // @[LoadQueue.scala 192:43:@35252.4]
  wire  _T_88428; // @[LoadQueue.scala 192:43:@35253.4]
  wire  _T_88429; // @[LoadQueue.scala 192:43:@35254.4]
  wire  _T_88430; // @[LoadQueue.scala 192:43:@35255.4]
  wire  _T_88431; // @[LoadQueue.scala 192:43:@35256.4]
  wire  _T_88432; // @[LoadQueue.scala 192:43:@35257.4]
  wire  _T_88433; // @[LoadQueue.scala 192:43:@35258.4]
  wire  _T_88434; // @[LoadQueue.scala 192:43:@35259.4]
  wire  _GEN_930; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_931; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_932; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_933; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_934; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_935; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_936; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_937; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_938; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_939; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_940; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_941; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_942; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_943; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_944; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_945; // @[LoadQueue.scala 193:43:@35261.6]
  wire  _GEN_947; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_948; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_949; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_950; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_951; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_952; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_953; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_954; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_955; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_956; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_957; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_958; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_959; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_960; // @[LoadQueue.scala 194:31:@35262.6]
  wire  _GEN_961; // @[LoadQueue.scala 194:31:@35262.6]
  wire [31:0] _GEN_963; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_964; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_965; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_966; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_967; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_968; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_969; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_970; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_971; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_972; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_973; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_974; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_975; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_976; // @[LoadQueue.scala 195:31:@35263.6]
  wire [31:0] _GEN_977; // @[LoadQueue.scala 195:31:@35263.6]
  wire  lastConflict_1_0; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_2; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_3; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_4; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_5; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_6; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_7; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_8; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_9; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_10; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_11; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_12; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_13; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_14; // @[LoadQueue.scala 192:53:@35260.4]
  wire  lastConflict_1_15; // @[LoadQueue.scala 192:53:@35260.4]
  wire  canBypass_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire [31:0] bypassVal_1; // @[LoadQueue.scala 192:53:@35260.4]
  wire [1:0] _T_88540; // @[LoadQueue.scala 191:60:@35317.4]
  wire [1:0] _T_88541; // @[LoadQueue.scala 191:60:@35318.4]
  wire [2:0] _T_88542; // @[LoadQueue.scala 191:60:@35319.4]
  wire [2:0] _T_88543; // @[LoadQueue.scala 191:60:@35320.4]
  wire [2:0] _T_88544; // @[LoadQueue.scala 191:60:@35321.4]
  wire [2:0] _T_88545; // @[LoadQueue.scala 191:60:@35322.4]
  wire [3:0] _T_88546; // @[LoadQueue.scala 191:60:@35323.4]
  wire [3:0] _T_88547; // @[LoadQueue.scala 191:60:@35324.4]
  wire [3:0] _T_88548; // @[LoadQueue.scala 191:60:@35325.4]
  wire [3:0] _T_88549; // @[LoadQueue.scala 191:60:@35326.4]
  wire [3:0] _T_88550; // @[LoadQueue.scala 191:60:@35327.4]
  wire [3:0] _T_88551; // @[LoadQueue.scala 191:60:@35328.4]
  wire [3:0] _T_88552; // @[LoadQueue.scala 191:60:@35329.4]
  wire [3:0] _T_88553; // @[LoadQueue.scala 191:60:@35330.4]
  wire  _T_88556; // @[LoadQueue.scala 192:43:@35332.4]
  wire  _T_88557; // @[LoadQueue.scala 192:43:@35333.4]
  wire  _T_88558; // @[LoadQueue.scala 192:43:@35334.4]
  wire  _T_88559; // @[LoadQueue.scala 192:43:@35335.4]
  wire  _T_88560; // @[LoadQueue.scala 192:43:@35336.4]
  wire  _T_88561; // @[LoadQueue.scala 192:43:@35337.4]
  wire  _T_88562; // @[LoadQueue.scala 192:43:@35338.4]
  wire  _T_88563; // @[LoadQueue.scala 192:43:@35339.4]
  wire  _T_88564; // @[LoadQueue.scala 192:43:@35340.4]
  wire  _T_88565; // @[LoadQueue.scala 192:43:@35341.4]
  wire  _T_88566; // @[LoadQueue.scala 192:43:@35342.4]
  wire  _T_88567; // @[LoadQueue.scala 192:43:@35343.4]
  wire  _T_88568; // @[LoadQueue.scala 192:43:@35344.4]
  wire  _T_88569; // @[LoadQueue.scala 192:43:@35345.4]
  wire  _T_88570; // @[LoadQueue.scala 192:43:@35346.4]
  wire  _GEN_996; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_997; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_998; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_999; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1000; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1001; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1002; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1003; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1004; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1005; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1006; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1007; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1008; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1009; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1010; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1011; // @[LoadQueue.scala 193:43:@35348.6]
  wire  _GEN_1013; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1014; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1015; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1016; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1017; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1018; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1019; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1020; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1021; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1022; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1023; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1024; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1025; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1026; // @[LoadQueue.scala 194:31:@35349.6]
  wire  _GEN_1027; // @[LoadQueue.scala 194:31:@35349.6]
  wire [31:0] _GEN_1029; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1030; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1031; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1032; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1033; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1034; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1035; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1036; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1037; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1038; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1039; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1040; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1041; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1042; // @[LoadQueue.scala 195:31:@35350.6]
  wire [31:0] _GEN_1043; // @[LoadQueue.scala 195:31:@35350.6]
  wire  lastConflict_2_0; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_1; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_3; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_4; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_5; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_6; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_7; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_8; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_9; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_10; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_11; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_12; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_13; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_14; // @[LoadQueue.scala 192:53:@35347.4]
  wire  lastConflict_2_15; // @[LoadQueue.scala 192:53:@35347.4]
  wire  canBypass_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire [31:0] bypassVal_2; // @[LoadQueue.scala 192:53:@35347.4]
  wire [1:0] _T_88676; // @[LoadQueue.scala 191:60:@35404.4]
  wire [1:0] _T_88677; // @[LoadQueue.scala 191:60:@35405.4]
  wire [2:0] _T_88678; // @[LoadQueue.scala 191:60:@35406.4]
  wire [2:0] _T_88679; // @[LoadQueue.scala 191:60:@35407.4]
  wire [2:0] _T_88680; // @[LoadQueue.scala 191:60:@35408.4]
  wire [2:0] _T_88681; // @[LoadQueue.scala 191:60:@35409.4]
  wire [3:0] _T_88682; // @[LoadQueue.scala 191:60:@35410.4]
  wire [3:0] _T_88683; // @[LoadQueue.scala 191:60:@35411.4]
  wire [3:0] _T_88684; // @[LoadQueue.scala 191:60:@35412.4]
  wire [3:0] _T_88685; // @[LoadQueue.scala 191:60:@35413.4]
  wire [3:0] _T_88686; // @[LoadQueue.scala 191:60:@35414.4]
  wire [3:0] _T_88687; // @[LoadQueue.scala 191:60:@35415.4]
  wire [3:0] _T_88688; // @[LoadQueue.scala 191:60:@35416.4]
  wire [3:0] _T_88689; // @[LoadQueue.scala 191:60:@35417.4]
  wire  _T_88692; // @[LoadQueue.scala 192:43:@35419.4]
  wire  _T_88693; // @[LoadQueue.scala 192:43:@35420.4]
  wire  _T_88694; // @[LoadQueue.scala 192:43:@35421.4]
  wire  _T_88695; // @[LoadQueue.scala 192:43:@35422.4]
  wire  _T_88696; // @[LoadQueue.scala 192:43:@35423.4]
  wire  _T_88697; // @[LoadQueue.scala 192:43:@35424.4]
  wire  _T_88698; // @[LoadQueue.scala 192:43:@35425.4]
  wire  _T_88699; // @[LoadQueue.scala 192:43:@35426.4]
  wire  _T_88700; // @[LoadQueue.scala 192:43:@35427.4]
  wire  _T_88701; // @[LoadQueue.scala 192:43:@35428.4]
  wire  _T_88702; // @[LoadQueue.scala 192:43:@35429.4]
  wire  _T_88703; // @[LoadQueue.scala 192:43:@35430.4]
  wire  _T_88704; // @[LoadQueue.scala 192:43:@35431.4]
  wire  _T_88705; // @[LoadQueue.scala 192:43:@35432.4]
  wire  _T_88706; // @[LoadQueue.scala 192:43:@35433.4]
  wire  _GEN_1062; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1063; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1064; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1065; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1066; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1067; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1068; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1069; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1070; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1071; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1072; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1073; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1074; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1075; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1076; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1077; // @[LoadQueue.scala 193:43:@35435.6]
  wire  _GEN_1079; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1080; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1081; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1082; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1083; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1084; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1085; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1086; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1087; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1088; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1089; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1090; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1091; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1092; // @[LoadQueue.scala 194:31:@35436.6]
  wire  _GEN_1093; // @[LoadQueue.scala 194:31:@35436.6]
  wire [31:0] _GEN_1095; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1096; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1097; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1098; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1099; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1100; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1101; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1102; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1103; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1104; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1105; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1106; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1107; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1108; // @[LoadQueue.scala 195:31:@35437.6]
  wire [31:0] _GEN_1109; // @[LoadQueue.scala 195:31:@35437.6]
  wire  lastConflict_3_0; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_1; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_2; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_4; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_5; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_6; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_7; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_8; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_9; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_10; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_11; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_12; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_13; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_14; // @[LoadQueue.scala 192:53:@35434.4]
  wire  lastConflict_3_15; // @[LoadQueue.scala 192:53:@35434.4]
  wire  canBypass_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire [31:0] bypassVal_3; // @[LoadQueue.scala 192:53:@35434.4]
  wire [1:0] _T_88812; // @[LoadQueue.scala 191:60:@35491.4]
  wire [1:0] _T_88813; // @[LoadQueue.scala 191:60:@35492.4]
  wire [2:0] _T_88814; // @[LoadQueue.scala 191:60:@35493.4]
  wire [2:0] _T_88815; // @[LoadQueue.scala 191:60:@35494.4]
  wire [2:0] _T_88816; // @[LoadQueue.scala 191:60:@35495.4]
  wire [2:0] _T_88817; // @[LoadQueue.scala 191:60:@35496.4]
  wire [3:0] _T_88818; // @[LoadQueue.scala 191:60:@35497.4]
  wire [3:0] _T_88819; // @[LoadQueue.scala 191:60:@35498.4]
  wire [3:0] _T_88820; // @[LoadQueue.scala 191:60:@35499.4]
  wire [3:0] _T_88821; // @[LoadQueue.scala 191:60:@35500.4]
  wire [3:0] _T_88822; // @[LoadQueue.scala 191:60:@35501.4]
  wire [3:0] _T_88823; // @[LoadQueue.scala 191:60:@35502.4]
  wire [3:0] _T_88824; // @[LoadQueue.scala 191:60:@35503.4]
  wire [3:0] _T_88825; // @[LoadQueue.scala 191:60:@35504.4]
  wire  _T_88828; // @[LoadQueue.scala 192:43:@35506.4]
  wire  _T_88829; // @[LoadQueue.scala 192:43:@35507.4]
  wire  _T_88830; // @[LoadQueue.scala 192:43:@35508.4]
  wire  _T_88831; // @[LoadQueue.scala 192:43:@35509.4]
  wire  _T_88832; // @[LoadQueue.scala 192:43:@35510.4]
  wire  _T_88833; // @[LoadQueue.scala 192:43:@35511.4]
  wire  _T_88834; // @[LoadQueue.scala 192:43:@35512.4]
  wire  _T_88835; // @[LoadQueue.scala 192:43:@35513.4]
  wire  _T_88836; // @[LoadQueue.scala 192:43:@35514.4]
  wire  _T_88837; // @[LoadQueue.scala 192:43:@35515.4]
  wire  _T_88838; // @[LoadQueue.scala 192:43:@35516.4]
  wire  _T_88839; // @[LoadQueue.scala 192:43:@35517.4]
  wire  _T_88840; // @[LoadQueue.scala 192:43:@35518.4]
  wire  _T_88841; // @[LoadQueue.scala 192:43:@35519.4]
  wire  _T_88842; // @[LoadQueue.scala 192:43:@35520.4]
  wire  _GEN_1128; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1129; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1130; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1131; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1132; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1133; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1134; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1135; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1136; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1137; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1138; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1139; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1140; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1141; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1142; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1143; // @[LoadQueue.scala 193:43:@35522.6]
  wire  _GEN_1145; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1146; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1147; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1148; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1149; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1150; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1151; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1152; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1153; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1154; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1155; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1156; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1157; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1158; // @[LoadQueue.scala 194:31:@35523.6]
  wire  _GEN_1159; // @[LoadQueue.scala 194:31:@35523.6]
  wire [31:0] _GEN_1161; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1162; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1163; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1164; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1165; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1166; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1167; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1168; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1169; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1170; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1171; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1172; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1173; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1174; // @[LoadQueue.scala 195:31:@35524.6]
  wire [31:0] _GEN_1175; // @[LoadQueue.scala 195:31:@35524.6]
  wire  lastConflict_4_0; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_1; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_2; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_3; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_5; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_6; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_7; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_8; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_9; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_10; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_11; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_12; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_13; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_14; // @[LoadQueue.scala 192:53:@35521.4]
  wire  lastConflict_4_15; // @[LoadQueue.scala 192:53:@35521.4]
  wire  canBypass_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire [31:0] bypassVal_4; // @[LoadQueue.scala 192:53:@35521.4]
  wire [1:0] _T_88948; // @[LoadQueue.scala 191:60:@35578.4]
  wire [1:0] _T_88949; // @[LoadQueue.scala 191:60:@35579.4]
  wire [2:0] _T_88950; // @[LoadQueue.scala 191:60:@35580.4]
  wire [2:0] _T_88951; // @[LoadQueue.scala 191:60:@35581.4]
  wire [2:0] _T_88952; // @[LoadQueue.scala 191:60:@35582.4]
  wire [2:0] _T_88953; // @[LoadQueue.scala 191:60:@35583.4]
  wire [3:0] _T_88954; // @[LoadQueue.scala 191:60:@35584.4]
  wire [3:0] _T_88955; // @[LoadQueue.scala 191:60:@35585.4]
  wire [3:0] _T_88956; // @[LoadQueue.scala 191:60:@35586.4]
  wire [3:0] _T_88957; // @[LoadQueue.scala 191:60:@35587.4]
  wire [3:0] _T_88958; // @[LoadQueue.scala 191:60:@35588.4]
  wire [3:0] _T_88959; // @[LoadQueue.scala 191:60:@35589.4]
  wire [3:0] _T_88960; // @[LoadQueue.scala 191:60:@35590.4]
  wire [3:0] _T_88961; // @[LoadQueue.scala 191:60:@35591.4]
  wire  _T_88964; // @[LoadQueue.scala 192:43:@35593.4]
  wire  _T_88965; // @[LoadQueue.scala 192:43:@35594.4]
  wire  _T_88966; // @[LoadQueue.scala 192:43:@35595.4]
  wire  _T_88967; // @[LoadQueue.scala 192:43:@35596.4]
  wire  _T_88968; // @[LoadQueue.scala 192:43:@35597.4]
  wire  _T_88969; // @[LoadQueue.scala 192:43:@35598.4]
  wire  _T_88970; // @[LoadQueue.scala 192:43:@35599.4]
  wire  _T_88971; // @[LoadQueue.scala 192:43:@35600.4]
  wire  _T_88972; // @[LoadQueue.scala 192:43:@35601.4]
  wire  _T_88973; // @[LoadQueue.scala 192:43:@35602.4]
  wire  _T_88974; // @[LoadQueue.scala 192:43:@35603.4]
  wire  _T_88975; // @[LoadQueue.scala 192:43:@35604.4]
  wire  _T_88976; // @[LoadQueue.scala 192:43:@35605.4]
  wire  _T_88977; // @[LoadQueue.scala 192:43:@35606.4]
  wire  _T_88978; // @[LoadQueue.scala 192:43:@35607.4]
  wire  _GEN_1194; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1195; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1196; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1197; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1198; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1199; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1200; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1201; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1202; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1203; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1204; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1205; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1206; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1207; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1208; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1209; // @[LoadQueue.scala 193:43:@35609.6]
  wire  _GEN_1211; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1212; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1213; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1214; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1215; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1216; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1217; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1218; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1219; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1220; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1221; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1222; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1223; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1224; // @[LoadQueue.scala 194:31:@35610.6]
  wire  _GEN_1225; // @[LoadQueue.scala 194:31:@35610.6]
  wire [31:0] _GEN_1227; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1228; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1229; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1230; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1231; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1232; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1233; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1234; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1235; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1236; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1237; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1238; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1239; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1240; // @[LoadQueue.scala 195:31:@35611.6]
  wire [31:0] _GEN_1241; // @[LoadQueue.scala 195:31:@35611.6]
  wire  lastConflict_5_0; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_1; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_2; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_3; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_4; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_6; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_7; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_8; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_9; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_10; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_11; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_12; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_13; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_14; // @[LoadQueue.scala 192:53:@35608.4]
  wire  lastConflict_5_15; // @[LoadQueue.scala 192:53:@35608.4]
  wire  canBypass_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire [31:0] bypassVal_5; // @[LoadQueue.scala 192:53:@35608.4]
  wire [1:0] _T_89084; // @[LoadQueue.scala 191:60:@35665.4]
  wire [1:0] _T_89085; // @[LoadQueue.scala 191:60:@35666.4]
  wire [2:0] _T_89086; // @[LoadQueue.scala 191:60:@35667.4]
  wire [2:0] _T_89087; // @[LoadQueue.scala 191:60:@35668.4]
  wire [2:0] _T_89088; // @[LoadQueue.scala 191:60:@35669.4]
  wire [2:0] _T_89089; // @[LoadQueue.scala 191:60:@35670.4]
  wire [3:0] _T_89090; // @[LoadQueue.scala 191:60:@35671.4]
  wire [3:0] _T_89091; // @[LoadQueue.scala 191:60:@35672.4]
  wire [3:0] _T_89092; // @[LoadQueue.scala 191:60:@35673.4]
  wire [3:0] _T_89093; // @[LoadQueue.scala 191:60:@35674.4]
  wire [3:0] _T_89094; // @[LoadQueue.scala 191:60:@35675.4]
  wire [3:0] _T_89095; // @[LoadQueue.scala 191:60:@35676.4]
  wire [3:0] _T_89096; // @[LoadQueue.scala 191:60:@35677.4]
  wire [3:0] _T_89097; // @[LoadQueue.scala 191:60:@35678.4]
  wire  _T_89100; // @[LoadQueue.scala 192:43:@35680.4]
  wire  _T_89101; // @[LoadQueue.scala 192:43:@35681.4]
  wire  _T_89102; // @[LoadQueue.scala 192:43:@35682.4]
  wire  _T_89103; // @[LoadQueue.scala 192:43:@35683.4]
  wire  _T_89104; // @[LoadQueue.scala 192:43:@35684.4]
  wire  _T_89105; // @[LoadQueue.scala 192:43:@35685.4]
  wire  _T_89106; // @[LoadQueue.scala 192:43:@35686.4]
  wire  _T_89107; // @[LoadQueue.scala 192:43:@35687.4]
  wire  _T_89108; // @[LoadQueue.scala 192:43:@35688.4]
  wire  _T_89109; // @[LoadQueue.scala 192:43:@35689.4]
  wire  _T_89110; // @[LoadQueue.scala 192:43:@35690.4]
  wire  _T_89111; // @[LoadQueue.scala 192:43:@35691.4]
  wire  _T_89112; // @[LoadQueue.scala 192:43:@35692.4]
  wire  _T_89113; // @[LoadQueue.scala 192:43:@35693.4]
  wire  _T_89114; // @[LoadQueue.scala 192:43:@35694.4]
  wire  _GEN_1260; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1261; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1262; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1263; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1264; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1265; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1266; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1267; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1268; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1269; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1270; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1271; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1272; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1273; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1274; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1275; // @[LoadQueue.scala 193:43:@35696.6]
  wire  _GEN_1277; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1278; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1279; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1280; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1281; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1282; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1283; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1284; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1285; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1286; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1287; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1288; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1289; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1290; // @[LoadQueue.scala 194:31:@35697.6]
  wire  _GEN_1291; // @[LoadQueue.scala 194:31:@35697.6]
  wire [31:0] _GEN_1293; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1294; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1295; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1296; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1297; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1298; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1299; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1300; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1301; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1302; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1303; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1304; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1305; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1306; // @[LoadQueue.scala 195:31:@35698.6]
  wire [31:0] _GEN_1307; // @[LoadQueue.scala 195:31:@35698.6]
  wire  lastConflict_6_0; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_1; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_2; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_3; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_4; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_5; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_7; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_8; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_9; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_10; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_11; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_12; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_13; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_14; // @[LoadQueue.scala 192:53:@35695.4]
  wire  lastConflict_6_15; // @[LoadQueue.scala 192:53:@35695.4]
  wire  canBypass_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire [31:0] bypassVal_6; // @[LoadQueue.scala 192:53:@35695.4]
  wire [1:0] _T_89220; // @[LoadQueue.scala 191:60:@35752.4]
  wire [1:0] _T_89221; // @[LoadQueue.scala 191:60:@35753.4]
  wire [2:0] _T_89222; // @[LoadQueue.scala 191:60:@35754.4]
  wire [2:0] _T_89223; // @[LoadQueue.scala 191:60:@35755.4]
  wire [2:0] _T_89224; // @[LoadQueue.scala 191:60:@35756.4]
  wire [2:0] _T_89225; // @[LoadQueue.scala 191:60:@35757.4]
  wire [3:0] _T_89226; // @[LoadQueue.scala 191:60:@35758.4]
  wire [3:0] _T_89227; // @[LoadQueue.scala 191:60:@35759.4]
  wire [3:0] _T_89228; // @[LoadQueue.scala 191:60:@35760.4]
  wire [3:0] _T_89229; // @[LoadQueue.scala 191:60:@35761.4]
  wire [3:0] _T_89230; // @[LoadQueue.scala 191:60:@35762.4]
  wire [3:0] _T_89231; // @[LoadQueue.scala 191:60:@35763.4]
  wire [3:0] _T_89232; // @[LoadQueue.scala 191:60:@35764.4]
  wire [3:0] _T_89233; // @[LoadQueue.scala 191:60:@35765.4]
  wire  _T_89236; // @[LoadQueue.scala 192:43:@35767.4]
  wire  _T_89237; // @[LoadQueue.scala 192:43:@35768.4]
  wire  _T_89238; // @[LoadQueue.scala 192:43:@35769.4]
  wire  _T_89239; // @[LoadQueue.scala 192:43:@35770.4]
  wire  _T_89240; // @[LoadQueue.scala 192:43:@35771.4]
  wire  _T_89241; // @[LoadQueue.scala 192:43:@35772.4]
  wire  _T_89242; // @[LoadQueue.scala 192:43:@35773.4]
  wire  _T_89243; // @[LoadQueue.scala 192:43:@35774.4]
  wire  _T_89244; // @[LoadQueue.scala 192:43:@35775.4]
  wire  _T_89245; // @[LoadQueue.scala 192:43:@35776.4]
  wire  _T_89246; // @[LoadQueue.scala 192:43:@35777.4]
  wire  _T_89247; // @[LoadQueue.scala 192:43:@35778.4]
  wire  _T_89248; // @[LoadQueue.scala 192:43:@35779.4]
  wire  _T_89249; // @[LoadQueue.scala 192:43:@35780.4]
  wire  _T_89250; // @[LoadQueue.scala 192:43:@35781.4]
  wire  _GEN_1326; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1327; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1328; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1329; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1330; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1331; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1332; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1333; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1334; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1335; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1336; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1337; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1338; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1339; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1340; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1341; // @[LoadQueue.scala 193:43:@35783.6]
  wire  _GEN_1343; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1344; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1345; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1346; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1347; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1348; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1349; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1350; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1351; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1352; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1353; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1354; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1355; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1356; // @[LoadQueue.scala 194:31:@35784.6]
  wire  _GEN_1357; // @[LoadQueue.scala 194:31:@35784.6]
  wire [31:0] _GEN_1359; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1360; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1361; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1362; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1363; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1364; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1365; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1366; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1367; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1368; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1369; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1370; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1371; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1372; // @[LoadQueue.scala 195:31:@35785.6]
  wire [31:0] _GEN_1373; // @[LoadQueue.scala 195:31:@35785.6]
  wire  lastConflict_7_0; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_1; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_2; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_3; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_4; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_5; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_6; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_8; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_9; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_10; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_11; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_12; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_13; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_14; // @[LoadQueue.scala 192:53:@35782.4]
  wire  lastConflict_7_15; // @[LoadQueue.scala 192:53:@35782.4]
  wire  canBypass_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire [31:0] bypassVal_7; // @[LoadQueue.scala 192:53:@35782.4]
  wire [1:0] _T_89356; // @[LoadQueue.scala 191:60:@35839.4]
  wire [1:0] _T_89357; // @[LoadQueue.scala 191:60:@35840.4]
  wire [2:0] _T_89358; // @[LoadQueue.scala 191:60:@35841.4]
  wire [2:0] _T_89359; // @[LoadQueue.scala 191:60:@35842.4]
  wire [2:0] _T_89360; // @[LoadQueue.scala 191:60:@35843.4]
  wire [2:0] _T_89361; // @[LoadQueue.scala 191:60:@35844.4]
  wire [3:0] _T_89362; // @[LoadQueue.scala 191:60:@35845.4]
  wire [3:0] _T_89363; // @[LoadQueue.scala 191:60:@35846.4]
  wire [3:0] _T_89364; // @[LoadQueue.scala 191:60:@35847.4]
  wire [3:0] _T_89365; // @[LoadQueue.scala 191:60:@35848.4]
  wire [3:0] _T_89366; // @[LoadQueue.scala 191:60:@35849.4]
  wire [3:0] _T_89367; // @[LoadQueue.scala 191:60:@35850.4]
  wire [3:0] _T_89368; // @[LoadQueue.scala 191:60:@35851.4]
  wire [3:0] _T_89369; // @[LoadQueue.scala 191:60:@35852.4]
  wire  _T_89372; // @[LoadQueue.scala 192:43:@35854.4]
  wire  _T_89373; // @[LoadQueue.scala 192:43:@35855.4]
  wire  _T_89374; // @[LoadQueue.scala 192:43:@35856.4]
  wire  _T_89375; // @[LoadQueue.scala 192:43:@35857.4]
  wire  _T_89376; // @[LoadQueue.scala 192:43:@35858.4]
  wire  _T_89377; // @[LoadQueue.scala 192:43:@35859.4]
  wire  _T_89378; // @[LoadQueue.scala 192:43:@35860.4]
  wire  _T_89379; // @[LoadQueue.scala 192:43:@35861.4]
  wire  _T_89380; // @[LoadQueue.scala 192:43:@35862.4]
  wire  _T_89381; // @[LoadQueue.scala 192:43:@35863.4]
  wire  _T_89382; // @[LoadQueue.scala 192:43:@35864.4]
  wire  _T_89383; // @[LoadQueue.scala 192:43:@35865.4]
  wire  _T_89384; // @[LoadQueue.scala 192:43:@35866.4]
  wire  _T_89385; // @[LoadQueue.scala 192:43:@35867.4]
  wire  _T_89386; // @[LoadQueue.scala 192:43:@35868.4]
  wire  _GEN_1392; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1393; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1394; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1395; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1396; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1397; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1398; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1399; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1400; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1401; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1402; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1403; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1404; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1405; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1406; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1407; // @[LoadQueue.scala 193:43:@35870.6]
  wire  _GEN_1409; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1410; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1411; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1412; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1413; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1414; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1415; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1416; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1417; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1418; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1419; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1420; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1421; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1422; // @[LoadQueue.scala 194:31:@35871.6]
  wire  _GEN_1423; // @[LoadQueue.scala 194:31:@35871.6]
  wire [31:0] _GEN_1425; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1426; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1427; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1428; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1429; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1430; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1431; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1432; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1433; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1434; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1435; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1436; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1437; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1438; // @[LoadQueue.scala 195:31:@35872.6]
  wire [31:0] _GEN_1439; // @[LoadQueue.scala 195:31:@35872.6]
  wire  lastConflict_8_0; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_1; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_2; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_3; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_4; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_5; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_6; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_7; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_9; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_10; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_11; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_12; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_13; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_14; // @[LoadQueue.scala 192:53:@35869.4]
  wire  lastConflict_8_15; // @[LoadQueue.scala 192:53:@35869.4]
  wire  canBypass_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire [31:0] bypassVal_8; // @[LoadQueue.scala 192:53:@35869.4]
  wire [1:0] _T_89492; // @[LoadQueue.scala 191:60:@35926.4]
  wire [1:0] _T_89493; // @[LoadQueue.scala 191:60:@35927.4]
  wire [2:0] _T_89494; // @[LoadQueue.scala 191:60:@35928.4]
  wire [2:0] _T_89495; // @[LoadQueue.scala 191:60:@35929.4]
  wire [2:0] _T_89496; // @[LoadQueue.scala 191:60:@35930.4]
  wire [2:0] _T_89497; // @[LoadQueue.scala 191:60:@35931.4]
  wire [3:0] _T_89498; // @[LoadQueue.scala 191:60:@35932.4]
  wire [3:0] _T_89499; // @[LoadQueue.scala 191:60:@35933.4]
  wire [3:0] _T_89500; // @[LoadQueue.scala 191:60:@35934.4]
  wire [3:0] _T_89501; // @[LoadQueue.scala 191:60:@35935.4]
  wire [3:0] _T_89502; // @[LoadQueue.scala 191:60:@35936.4]
  wire [3:0] _T_89503; // @[LoadQueue.scala 191:60:@35937.4]
  wire [3:0] _T_89504; // @[LoadQueue.scala 191:60:@35938.4]
  wire [3:0] _T_89505; // @[LoadQueue.scala 191:60:@35939.4]
  wire  _T_89508; // @[LoadQueue.scala 192:43:@35941.4]
  wire  _T_89509; // @[LoadQueue.scala 192:43:@35942.4]
  wire  _T_89510; // @[LoadQueue.scala 192:43:@35943.4]
  wire  _T_89511; // @[LoadQueue.scala 192:43:@35944.4]
  wire  _T_89512; // @[LoadQueue.scala 192:43:@35945.4]
  wire  _T_89513; // @[LoadQueue.scala 192:43:@35946.4]
  wire  _T_89514; // @[LoadQueue.scala 192:43:@35947.4]
  wire  _T_89515; // @[LoadQueue.scala 192:43:@35948.4]
  wire  _T_89516; // @[LoadQueue.scala 192:43:@35949.4]
  wire  _T_89517; // @[LoadQueue.scala 192:43:@35950.4]
  wire  _T_89518; // @[LoadQueue.scala 192:43:@35951.4]
  wire  _T_89519; // @[LoadQueue.scala 192:43:@35952.4]
  wire  _T_89520; // @[LoadQueue.scala 192:43:@35953.4]
  wire  _T_89521; // @[LoadQueue.scala 192:43:@35954.4]
  wire  _T_89522; // @[LoadQueue.scala 192:43:@35955.4]
  wire  _GEN_1458; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1459; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1460; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1461; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1462; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1463; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1464; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1465; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1466; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1467; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1468; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1469; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1470; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1471; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1472; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1473; // @[LoadQueue.scala 193:43:@35957.6]
  wire  _GEN_1475; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1476; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1477; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1478; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1479; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1480; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1481; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1482; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1483; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1484; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1485; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1486; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1487; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1488; // @[LoadQueue.scala 194:31:@35958.6]
  wire  _GEN_1489; // @[LoadQueue.scala 194:31:@35958.6]
  wire [31:0] _GEN_1491; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1492; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1493; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1494; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1495; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1496; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1497; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1498; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1499; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1500; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1501; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1502; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1503; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1504; // @[LoadQueue.scala 195:31:@35959.6]
  wire [31:0] _GEN_1505; // @[LoadQueue.scala 195:31:@35959.6]
  wire  lastConflict_9_0; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_1; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_2; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_3; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_4; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_5; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_6; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_7; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_8; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_10; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_11; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_12; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_13; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_14; // @[LoadQueue.scala 192:53:@35956.4]
  wire  lastConflict_9_15; // @[LoadQueue.scala 192:53:@35956.4]
  wire  canBypass_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire [31:0] bypassVal_9; // @[LoadQueue.scala 192:53:@35956.4]
  wire [1:0] _T_89628; // @[LoadQueue.scala 191:60:@36013.4]
  wire [1:0] _T_89629; // @[LoadQueue.scala 191:60:@36014.4]
  wire [2:0] _T_89630; // @[LoadQueue.scala 191:60:@36015.4]
  wire [2:0] _T_89631; // @[LoadQueue.scala 191:60:@36016.4]
  wire [2:0] _T_89632; // @[LoadQueue.scala 191:60:@36017.4]
  wire [2:0] _T_89633; // @[LoadQueue.scala 191:60:@36018.4]
  wire [3:0] _T_89634; // @[LoadQueue.scala 191:60:@36019.4]
  wire [3:0] _T_89635; // @[LoadQueue.scala 191:60:@36020.4]
  wire [3:0] _T_89636; // @[LoadQueue.scala 191:60:@36021.4]
  wire [3:0] _T_89637; // @[LoadQueue.scala 191:60:@36022.4]
  wire [3:0] _T_89638; // @[LoadQueue.scala 191:60:@36023.4]
  wire [3:0] _T_89639; // @[LoadQueue.scala 191:60:@36024.4]
  wire [3:0] _T_89640; // @[LoadQueue.scala 191:60:@36025.4]
  wire [3:0] _T_89641; // @[LoadQueue.scala 191:60:@36026.4]
  wire  _T_89644; // @[LoadQueue.scala 192:43:@36028.4]
  wire  _T_89645; // @[LoadQueue.scala 192:43:@36029.4]
  wire  _T_89646; // @[LoadQueue.scala 192:43:@36030.4]
  wire  _T_89647; // @[LoadQueue.scala 192:43:@36031.4]
  wire  _T_89648; // @[LoadQueue.scala 192:43:@36032.4]
  wire  _T_89649; // @[LoadQueue.scala 192:43:@36033.4]
  wire  _T_89650; // @[LoadQueue.scala 192:43:@36034.4]
  wire  _T_89651; // @[LoadQueue.scala 192:43:@36035.4]
  wire  _T_89652; // @[LoadQueue.scala 192:43:@36036.4]
  wire  _T_89653; // @[LoadQueue.scala 192:43:@36037.4]
  wire  _T_89654; // @[LoadQueue.scala 192:43:@36038.4]
  wire  _T_89655; // @[LoadQueue.scala 192:43:@36039.4]
  wire  _T_89656; // @[LoadQueue.scala 192:43:@36040.4]
  wire  _T_89657; // @[LoadQueue.scala 192:43:@36041.4]
  wire  _T_89658; // @[LoadQueue.scala 192:43:@36042.4]
  wire  _GEN_1524; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1525; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1526; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1527; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1528; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1529; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1530; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1531; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1532; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1533; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1534; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1535; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1536; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1537; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1538; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1539; // @[LoadQueue.scala 193:43:@36044.6]
  wire  _GEN_1541; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1542; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1543; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1544; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1545; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1546; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1547; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1548; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1549; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1550; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1551; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1552; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1553; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1554; // @[LoadQueue.scala 194:31:@36045.6]
  wire  _GEN_1555; // @[LoadQueue.scala 194:31:@36045.6]
  wire [31:0] _GEN_1557; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1558; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1559; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1560; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1561; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1562; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1563; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1564; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1565; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1566; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1567; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1568; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1569; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1570; // @[LoadQueue.scala 195:31:@36046.6]
  wire [31:0] _GEN_1571; // @[LoadQueue.scala 195:31:@36046.6]
  wire  lastConflict_10_0; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_1; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_2; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_3; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_4; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_5; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_6; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_7; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_8; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_9; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_11; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_12; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_13; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_14; // @[LoadQueue.scala 192:53:@36043.4]
  wire  lastConflict_10_15; // @[LoadQueue.scala 192:53:@36043.4]
  wire  canBypass_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire [31:0] bypassVal_10; // @[LoadQueue.scala 192:53:@36043.4]
  wire [1:0] _T_89764; // @[LoadQueue.scala 191:60:@36100.4]
  wire [1:0] _T_89765; // @[LoadQueue.scala 191:60:@36101.4]
  wire [2:0] _T_89766; // @[LoadQueue.scala 191:60:@36102.4]
  wire [2:0] _T_89767; // @[LoadQueue.scala 191:60:@36103.4]
  wire [2:0] _T_89768; // @[LoadQueue.scala 191:60:@36104.4]
  wire [2:0] _T_89769; // @[LoadQueue.scala 191:60:@36105.4]
  wire [3:0] _T_89770; // @[LoadQueue.scala 191:60:@36106.4]
  wire [3:0] _T_89771; // @[LoadQueue.scala 191:60:@36107.4]
  wire [3:0] _T_89772; // @[LoadQueue.scala 191:60:@36108.4]
  wire [3:0] _T_89773; // @[LoadQueue.scala 191:60:@36109.4]
  wire [3:0] _T_89774; // @[LoadQueue.scala 191:60:@36110.4]
  wire [3:0] _T_89775; // @[LoadQueue.scala 191:60:@36111.4]
  wire [3:0] _T_89776; // @[LoadQueue.scala 191:60:@36112.4]
  wire [3:0] _T_89777; // @[LoadQueue.scala 191:60:@36113.4]
  wire  _T_89780; // @[LoadQueue.scala 192:43:@36115.4]
  wire  _T_89781; // @[LoadQueue.scala 192:43:@36116.4]
  wire  _T_89782; // @[LoadQueue.scala 192:43:@36117.4]
  wire  _T_89783; // @[LoadQueue.scala 192:43:@36118.4]
  wire  _T_89784; // @[LoadQueue.scala 192:43:@36119.4]
  wire  _T_89785; // @[LoadQueue.scala 192:43:@36120.4]
  wire  _T_89786; // @[LoadQueue.scala 192:43:@36121.4]
  wire  _T_89787; // @[LoadQueue.scala 192:43:@36122.4]
  wire  _T_89788; // @[LoadQueue.scala 192:43:@36123.4]
  wire  _T_89789; // @[LoadQueue.scala 192:43:@36124.4]
  wire  _T_89790; // @[LoadQueue.scala 192:43:@36125.4]
  wire  _T_89791; // @[LoadQueue.scala 192:43:@36126.4]
  wire  _T_89792; // @[LoadQueue.scala 192:43:@36127.4]
  wire  _T_89793; // @[LoadQueue.scala 192:43:@36128.4]
  wire  _T_89794; // @[LoadQueue.scala 192:43:@36129.4]
  wire  _GEN_1590; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1591; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1592; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1593; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1594; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1595; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1596; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1597; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1598; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1599; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1600; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1601; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1602; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1603; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1604; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1605; // @[LoadQueue.scala 193:43:@36131.6]
  wire  _GEN_1607; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1608; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1609; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1610; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1611; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1612; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1613; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1614; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1615; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1616; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1617; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1618; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1619; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1620; // @[LoadQueue.scala 194:31:@36132.6]
  wire  _GEN_1621; // @[LoadQueue.scala 194:31:@36132.6]
  wire [31:0] _GEN_1623; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1624; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1625; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1626; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1627; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1628; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1629; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1630; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1631; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1632; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1633; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1634; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1635; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1636; // @[LoadQueue.scala 195:31:@36133.6]
  wire [31:0] _GEN_1637; // @[LoadQueue.scala 195:31:@36133.6]
  wire  lastConflict_11_0; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_1; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_2; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_3; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_4; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_5; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_6; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_7; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_8; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_9; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_10; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_12; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_13; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_14; // @[LoadQueue.scala 192:53:@36130.4]
  wire  lastConflict_11_15; // @[LoadQueue.scala 192:53:@36130.4]
  wire  canBypass_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire [31:0] bypassVal_11; // @[LoadQueue.scala 192:53:@36130.4]
  wire [1:0] _T_89900; // @[LoadQueue.scala 191:60:@36187.4]
  wire [1:0] _T_89901; // @[LoadQueue.scala 191:60:@36188.4]
  wire [2:0] _T_89902; // @[LoadQueue.scala 191:60:@36189.4]
  wire [2:0] _T_89903; // @[LoadQueue.scala 191:60:@36190.4]
  wire [2:0] _T_89904; // @[LoadQueue.scala 191:60:@36191.4]
  wire [2:0] _T_89905; // @[LoadQueue.scala 191:60:@36192.4]
  wire [3:0] _T_89906; // @[LoadQueue.scala 191:60:@36193.4]
  wire [3:0] _T_89907; // @[LoadQueue.scala 191:60:@36194.4]
  wire [3:0] _T_89908; // @[LoadQueue.scala 191:60:@36195.4]
  wire [3:0] _T_89909; // @[LoadQueue.scala 191:60:@36196.4]
  wire [3:0] _T_89910; // @[LoadQueue.scala 191:60:@36197.4]
  wire [3:0] _T_89911; // @[LoadQueue.scala 191:60:@36198.4]
  wire [3:0] _T_89912; // @[LoadQueue.scala 191:60:@36199.4]
  wire [3:0] _T_89913; // @[LoadQueue.scala 191:60:@36200.4]
  wire  _T_89916; // @[LoadQueue.scala 192:43:@36202.4]
  wire  _T_89917; // @[LoadQueue.scala 192:43:@36203.4]
  wire  _T_89918; // @[LoadQueue.scala 192:43:@36204.4]
  wire  _T_89919; // @[LoadQueue.scala 192:43:@36205.4]
  wire  _T_89920; // @[LoadQueue.scala 192:43:@36206.4]
  wire  _T_89921; // @[LoadQueue.scala 192:43:@36207.4]
  wire  _T_89922; // @[LoadQueue.scala 192:43:@36208.4]
  wire  _T_89923; // @[LoadQueue.scala 192:43:@36209.4]
  wire  _T_89924; // @[LoadQueue.scala 192:43:@36210.4]
  wire  _T_89925; // @[LoadQueue.scala 192:43:@36211.4]
  wire  _T_89926; // @[LoadQueue.scala 192:43:@36212.4]
  wire  _T_89927; // @[LoadQueue.scala 192:43:@36213.4]
  wire  _T_89928; // @[LoadQueue.scala 192:43:@36214.4]
  wire  _T_89929; // @[LoadQueue.scala 192:43:@36215.4]
  wire  _T_89930; // @[LoadQueue.scala 192:43:@36216.4]
  wire  _GEN_1656; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1657; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1658; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1659; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1660; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1661; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1662; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1663; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1664; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1665; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1666; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1667; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1668; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1669; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1670; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1671; // @[LoadQueue.scala 193:43:@36218.6]
  wire  _GEN_1673; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1674; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1675; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1676; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1677; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1678; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1679; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1680; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1681; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1682; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1683; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1684; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1685; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1686; // @[LoadQueue.scala 194:31:@36219.6]
  wire  _GEN_1687; // @[LoadQueue.scala 194:31:@36219.6]
  wire [31:0] _GEN_1689; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1690; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1691; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1692; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1693; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1694; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1695; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1696; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1697; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1698; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1699; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1700; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1701; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1702; // @[LoadQueue.scala 195:31:@36220.6]
  wire [31:0] _GEN_1703; // @[LoadQueue.scala 195:31:@36220.6]
  wire  lastConflict_12_0; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_1; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_2; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_3; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_4; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_5; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_6; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_7; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_8; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_9; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_10; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_11; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_13; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_14; // @[LoadQueue.scala 192:53:@36217.4]
  wire  lastConflict_12_15; // @[LoadQueue.scala 192:53:@36217.4]
  wire  canBypass_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire [31:0] bypassVal_12; // @[LoadQueue.scala 192:53:@36217.4]
  wire [1:0] _T_90036; // @[LoadQueue.scala 191:60:@36274.4]
  wire [1:0] _T_90037; // @[LoadQueue.scala 191:60:@36275.4]
  wire [2:0] _T_90038; // @[LoadQueue.scala 191:60:@36276.4]
  wire [2:0] _T_90039; // @[LoadQueue.scala 191:60:@36277.4]
  wire [2:0] _T_90040; // @[LoadQueue.scala 191:60:@36278.4]
  wire [2:0] _T_90041; // @[LoadQueue.scala 191:60:@36279.4]
  wire [3:0] _T_90042; // @[LoadQueue.scala 191:60:@36280.4]
  wire [3:0] _T_90043; // @[LoadQueue.scala 191:60:@36281.4]
  wire [3:0] _T_90044; // @[LoadQueue.scala 191:60:@36282.4]
  wire [3:0] _T_90045; // @[LoadQueue.scala 191:60:@36283.4]
  wire [3:0] _T_90046; // @[LoadQueue.scala 191:60:@36284.4]
  wire [3:0] _T_90047; // @[LoadQueue.scala 191:60:@36285.4]
  wire [3:0] _T_90048; // @[LoadQueue.scala 191:60:@36286.4]
  wire [3:0] _T_90049; // @[LoadQueue.scala 191:60:@36287.4]
  wire  _T_90052; // @[LoadQueue.scala 192:43:@36289.4]
  wire  _T_90053; // @[LoadQueue.scala 192:43:@36290.4]
  wire  _T_90054; // @[LoadQueue.scala 192:43:@36291.4]
  wire  _T_90055; // @[LoadQueue.scala 192:43:@36292.4]
  wire  _T_90056; // @[LoadQueue.scala 192:43:@36293.4]
  wire  _T_90057; // @[LoadQueue.scala 192:43:@36294.4]
  wire  _T_90058; // @[LoadQueue.scala 192:43:@36295.4]
  wire  _T_90059; // @[LoadQueue.scala 192:43:@36296.4]
  wire  _T_90060; // @[LoadQueue.scala 192:43:@36297.4]
  wire  _T_90061; // @[LoadQueue.scala 192:43:@36298.4]
  wire  _T_90062; // @[LoadQueue.scala 192:43:@36299.4]
  wire  _T_90063; // @[LoadQueue.scala 192:43:@36300.4]
  wire  _T_90064; // @[LoadQueue.scala 192:43:@36301.4]
  wire  _T_90065; // @[LoadQueue.scala 192:43:@36302.4]
  wire  _T_90066; // @[LoadQueue.scala 192:43:@36303.4]
  wire  _GEN_1722; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1723; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1724; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1725; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1726; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1727; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1728; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1729; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1730; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1731; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1732; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1733; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1734; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1735; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1736; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1737; // @[LoadQueue.scala 193:43:@36305.6]
  wire  _GEN_1739; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1740; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1741; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1742; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1743; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1744; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1745; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1746; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1747; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1748; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1749; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1750; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1751; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1752; // @[LoadQueue.scala 194:31:@36306.6]
  wire  _GEN_1753; // @[LoadQueue.scala 194:31:@36306.6]
  wire [31:0] _GEN_1755; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1756; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1757; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1758; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1759; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1760; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1761; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1762; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1763; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1764; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1765; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1766; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1767; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1768; // @[LoadQueue.scala 195:31:@36307.6]
  wire [31:0] _GEN_1769; // @[LoadQueue.scala 195:31:@36307.6]
  wire  lastConflict_13_0; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_1; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_2; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_3; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_4; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_5; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_6; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_7; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_8; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_9; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_10; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_11; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_12; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_14; // @[LoadQueue.scala 192:53:@36304.4]
  wire  lastConflict_13_15; // @[LoadQueue.scala 192:53:@36304.4]
  wire  canBypass_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire [31:0] bypassVal_13; // @[LoadQueue.scala 192:53:@36304.4]
  wire [1:0] _T_90172; // @[LoadQueue.scala 191:60:@36361.4]
  wire [1:0] _T_90173; // @[LoadQueue.scala 191:60:@36362.4]
  wire [2:0] _T_90174; // @[LoadQueue.scala 191:60:@36363.4]
  wire [2:0] _T_90175; // @[LoadQueue.scala 191:60:@36364.4]
  wire [2:0] _T_90176; // @[LoadQueue.scala 191:60:@36365.4]
  wire [2:0] _T_90177; // @[LoadQueue.scala 191:60:@36366.4]
  wire [3:0] _T_90178; // @[LoadQueue.scala 191:60:@36367.4]
  wire [3:0] _T_90179; // @[LoadQueue.scala 191:60:@36368.4]
  wire [3:0] _T_90180; // @[LoadQueue.scala 191:60:@36369.4]
  wire [3:0] _T_90181; // @[LoadQueue.scala 191:60:@36370.4]
  wire [3:0] _T_90182; // @[LoadQueue.scala 191:60:@36371.4]
  wire [3:0] _T_90183; // @[LoadQueue.scala 191:60:@36372.4]
  wire [3:0] _T_90184; // @[LoadQueue.scala 191:60:@36373.4]
  wire [3:0] _T_90185; // @[LoadQueue.scala 191:60:@36374.4]
  wire  _T_90188; // @[LoadQueue.scala 192:43:@36376.4]
  wire  _T_90189; // @[LoadQueue.scala 192:43:@36377.4]
  wire  _T_90190; // @[LoadQueue.scala 192:43:@36378.4]
  wire  _T_90191; // @[LoadQueue.scala 192:43:@36379.4]
  wire  _T_90192; // @[LoadQueue.scala 192:43:@36380.4]
  wire  _T_90193; // @[LoadQueue.scala 192:43:@36381.4]
  wire  _T_90194; // @[LoadQueue.scala 192:43:@36382.4]
  wire  _T_90195; // @[LoadQueue.scala 192:43:@36383.4]
  wire  _T_90196; // @[LoadQueue.scala 192:43:@36384.4]
  wire  _T_90197; // @[LoadQueue.scala 192:43:@36385.4]
  wire  _T_90198; // @[LoadQueue.scala 192:43:@36386.4]
  wire  _T_90199; // @[LoadQueue.scala 192:43:@36387.4]
  wire  _T_90200; // @[LoadQueue.scala 192:43:@36388.4]
  wire  _T_90201; // @[LoadQueue.scala 192:43:@36389.4]
  wire  _T_90202; // @[LoadQueue.scala 192:43:@36390.4]
  wire  _GEN_1788; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1789; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1790; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1791; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1792; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1793; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1794; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1795; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1796; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1797; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1798; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1799; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1800; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1801; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1802; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1803; // @[LoadQueue.scala 193:43:@36392.6]
  wire  _GEN_1805; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1806; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1807; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1808; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1809; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1810; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1811; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1812; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1813; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1814; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1815; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1816; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1817; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1818; // @[LoadQueue.scala 194:31:@36393.6]
  wire  _GEN_1819; // @[LoadQueue.scala 194:31:@36393.6]
  wire [31:0] _GEN_1821; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1822; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1823; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1824; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1825; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1826; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1827; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1828; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1829; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1830; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1831; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1832; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1833; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1834; // @[LoadQueue.scala 195:31:@36394.6]
  wire [31:0] _GEN_1835; // @[LoadQueue.scala 195:31:@36394.6]
  wire  lastConflict_14_0; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_1; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_2; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_3; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_4; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_5; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_6; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_7; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_8; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_9; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_10; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_11; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_12; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_13; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire  lastConflict_14_15; // @[LoadQueue.scala 192:53:@36391.4]
  wire  canBypass_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire [31:0] bypassVal_14; // @[LoadQueue.scala 192:53:@36391.4]
  wire [1:0] _T_90308; // @[LoadQueue.scala 191:60:@36448.4]
  wire [1:0] _T_90309; // @[LoadQueue.scala 191:60:@36449.4]
  wire [2:0] _T_90310; // @[LoadQueue.scala 191:60:@36450.4]
  wire [2:0] _T_90311; // @[LoadQueue.scala 191:60:@36451.4]
  wire [2:0] _T_90312; // @[LoadQueue.scala 191:60:@36452.4]
  wire [2:0] _T_90313; // @[LoadQueue.scala 191:60:@36453.4]
  wire [3:0] _T_90314; // @[LoadQueue.scala 191:60:@36454.4]
  wire [3:0] _T_90315; // @[LoadQueue.scala 191:60:@36455.4]
  wire [3:0] _T_90316; // @[LoadQueue.scala 191:60:@36456.4]
  wire [3:0] _T_90317; // @[LoadQueue.scala 191:60:@36457.4]
  wire [3:0] _T_90318; // @[LoadQueue.scala 191:60:@36458.4]
  wire [3:0] _T_90319; // @[LoadQueue.scala 191:60:@36459.4]
  wire [3:0] _T_90320; // @[LoadQueue.scala 191:60:@36460.4]
  wire [3:0] _T_90321; // @[LoadQueue.scala 191:60:@36461.4]
  wire  _T_90324; // @[LoadQueue.scala 192:43:@36463.4]
  wire  _T_90325; // @[LoadQueue.scala 192:43:@36464.4]
  wire  _T_90326; // @[LoadQueue.scala 192:43:@36465.4]
  wire  _T_90327; // @[LoadQueue.scala 192:43:@36466.4]
  wire  _T_90328; // @[LoadQueue.scala 192:43:@36467.4]
  wire  _T_90329; // @[LoadQueue.scala 192:43:@36468.4]
  wire  _T_90330; // @[LoadQueue.scala 192:43:@36469.4]
  wire  _T_90331; // @[LoadQueue.scala 192:43:@36470.4]
  wire  _T_90332; // @[LoadQueue.scala 192:43:@36471.4]
  wire  _T_90333; // @[LoadQueue.scala 192:43:@36472.4]
  wire  _T_90334; // @[LoadQueue.scala 192:43:@36473.4]
  wire  _T_90335; // @[LoadQueue.scala 192:43:@36474.4]
  wire  _T_90336; // @[LoadQueue.scala 192:43:@36475.4]
  wire  _T_90337; // @[LoadQueue.scala 192:43:@36476.4]
  wire  _T_90338; // @[LoadQueue.scala 192:43:@36477.4]
  wire  _GEN_1854; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1855; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1856; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1857; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1858; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1859; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1860; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1861; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1862; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1863; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1864; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1865; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1866; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1867; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1868; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1869; // @[LoadQueue.scala 193:43:@36479.6]
  wire  _GEN_1871; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1872; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1873; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1874; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1875; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1876; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1877; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1878; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1879; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1880; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1881; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1882; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1883; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1884; // @[LoadQueue.scala 194:31:@36480.6]
  wire  _GEN_1885; // @[LoadQueue.scala 194:31:@36480.6]
  wire [31:0] _GEN_1887; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1888; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1889; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1890; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1891; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1892; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1893; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1894; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1895; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1896; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1897; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1898; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1899; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1900; // @[LoadQueue.scala 195:31:@36481.6]
  wire [31:0] _GEN_1901; // @[LoadQueue.scala 195:31:@36481.6]
  wire  lastConflict_15_0; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_1; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_2; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_3; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_4; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_5; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_6; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_7; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_8; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_9; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_10; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_11; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_12; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_13; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_14; // @[LoadQueue.scala 192:53:@36478.4]
  wire  lastConflict_15_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire  canBypass_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire [31:0] bypassVal_15; // @[LoadQueue.scala 192:53:@36478.4]
  wire [15:0] _T_90398; // @[OneHot.scala 52:12:@36486.4]
  wire  _T_90400; // @[util.scala 33:60:@36488.4]
  wire  _T_90401; // @[util.scala 33:60:@36489.4]
  wire  _T_90402; // @[util.scala 33:60:@36490.4]
  wire  _T_90403; // @[util.scala 33:60:@36491.4]
  wire  _T_90404; // @[util.scala 33:60:@36492.4]
  wire  _T_90405; // @[util.scala 33:60:@36493.4]
  wire  _T_90406; // @[util.scala 33:60:@36494.4]
  wire  _T_90407; // @[util.scala 33:60:@36495.4]
  wire  _T_90408; // @[util.scala 33:60:@36496.4]
  wire  _T_90409; // @[util.scala 33:60:@36497.4]
  wire  _T_90410; // @[util.scala 33:60:@36498.4]
  wire  _T_90411; // @[util.scala 33:60:@36499.4]
  wire  _T_90412; // @[util.scala 33:60:@36500.4]
  wire  _T_90413; // @[util.scala 33:60:@36501.4]
  wire  _T_90414; // @[util.scala 33:60:@36502.4]
  wire  _T_90415; // @[util.scala 33:60:@36503.4]
  wire  _T_93512; // @[LoadQueue.scala 229:41:@39026.4]
  wire  _T_93513; // @[LoadQueue.scala 229:38:@39027.4]
  wire  _T_93515; // @[LoadQueue.scala 230:12:@39029.6]
  reg  prevPriorityRequest_15; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_739;
  wire  _T_93517; // @[LoadQueue.scala 230:46:@39030.6]
  wire  _T_93518; // @[LoadQueue.scala 230:43:@39031.6]
  wire  _T_93520; // @[LoadQueue.scala 230:84:@39032.6]
  wire  _T_93521; // @[LoadQueue.scala 230:81:@39033.6]
  wire  _T_93524; // @[LoadQueue.scala 233:86:@39036.8]
  wire  _T_93525; // @[LoadQueue.scala 233:86:@39037.8]
  wire  _T_93526; // @[LoadQueue.scala 233:86:@39038.8]
  wire  _T_93527; // @[LoadQueue.scala 233:86:@39039.8]
  wire  _T_93528; // @[LoadQueue.scala 233:86:@39040.8]
  wire  _T_93529; // @[LoadQueue.scala 233:86:@39041.8]
  wire  _T_93530; // @[LoadQueue.scala 233:86:@39042.8]
  wire  _T_93531; // @[LoadQueue.scala 233:86:@39043.8]
  wire  _T_93532; // @[LoadQueue.scala 233:86:@39044.8]
  wire  _T_93533; // @[LoadQueue.scala 233:86:@39045.8]
  wire  _T_93534; // @[LoadQueue.scala 233:86:@39046.8]
  wire  _T_93535; // @[LoadQueue.scala 233:86:@39047.8]
  wire  _T_93536; // @[LoadQueue.scala 233:86:@39048.8]
  wire  _T_93537; // @[LoadQueue.scala 233:86:@39049.8]
  wire  _T_93538; // @[LoadQueue.scala 233:86:@39050.8]
  wire  _T_93540; // @[LoadQueue.scala 233:38:@39051.8]
  wire  _T_93559; // @[LoadQueue.scala 234:11:@39068.8]
  wire  _T_93560; // @[LoadQueue.scala 233:103:@39069.8]
  wire  _GEN_2028; // @[LoadQueue.scala 230:110:@39034.6]
  wire  loadRequest_15; // @[LoadQueue.scala 229:71:@39028.4]
  wire [15:0] _T_90456; // @[Mux.scala 31:69:@36521.4]
  wire  _T_93428; // @[LoadQueue.scala 229:41:@38944.4]
  wire  _T_93429; // @[LoadQueue.scala 229:38:@38945.4]
  wire  _T_93431; // @[LoadQueue.scala 230:12:@38947.6]
  reg  prevPriorityRequest_14; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_740;
  wire  _T_93433; // @[LoadQueue.scala 230:46:@38948.6]
  wire  _T_93434; // @[LoadQueue.scala 230:43:@38949.6]
  wire  _T_93436; // @[LoadQueue.scala 230:84:@38950.6]
  wire  _T_93437; // @[LoadQueue.scala 230:81:@38951.6]
  wire  _T_93440; // @[LoadQueue.scala 233:86:@38954.8]
  wire  _T_93441; // @[LoadQueue.scala 233:86:@38955.8]
  wire  _T_93442; // @[LoadQueue.scala 233:86:@38956.8]
  wire  _T_93443; // @[LoadQueue.scala 233:86:@38957.8]
  wire  _T_93444; // @[LoadQueue.scala 233:86:@38958.8]
  wire  _T_93445; // @[LoadQueue.scala 233:86:@38959.8]
  wire  _T_93446; // @[LoadQueue.scala 233:86:@38960.8]
  wire  _T_93447; // @[LoadQueue.scala 233:86:@38961.8]
  wire  _T_93448; // @[LoadQueue.scala 233:86:@38962.8]
  wire  _T_93449; // @[LoadQueue.scala 233:86:@38963.8]
  wire  _T_93450; // @[LoadQueue.scala 233:86:@38964.8]
  wire  _T_93451; // @[LoadQueue.scala 233:86:@38965.8]
  wire  _T_93452; // @[LoadQueue.scala 233:86:@38966.8]
  wire  _T_93453; // @[LoadQueue.scala 233:86:@38967.8]
  wire  _T_93454; // @[LoadQueue.scala 233:86:@38968.8]
  wire  _T_93456; // @[LoadQueue.scala 233:38:@38969.8]
  wire  _T_93475; // @[LoadQueue.scala 234:11:@38986.8]
  wire  _T_93476; // @[LoadQueue.scala 233:103:@38987.8]
  wire  _GEN_2024; // @[LoadQueue.scala 230:110:@38952.6]
  wire  loadRequest_14; // @[LoadQueue.scala 229:71:@38946.4]
  wire [15:0] _T_90457; // @[Mux.scala 31:69:@36522.4]
  wire  _T_93344; // @[LoadQueue.scala 229:41:@38862.4]
  wire  _T_93345; // @[LoadQueue.scala 229:38:@38863.4]
  wire  _T_93347; // @[LoadQueue.scala 230:12:@38865.6]
  reg  prevPriorityRequest_13; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_741;
  wire  _T_93349; // @[LoadQueue.scala 230:46:@38866.6]
  wire  _T_93350; // @[LoadQueue.scala 230:43:@38867.6]
  wire  _T_93352; // @[LoadQueue.scala 230:84:@38868.6]
  wire  _T_93353; // @[LoadQueue.scala 230:81:@38869.6]
  wire  _T_93356; // @[LoadQueue.scala 233:86:@38872.8]
  wire  _T_93357; // @[LoadQueue.scala 233:86:@38873.8]
  wire  _T_93358; // @[LoadQueue.scala 233:86:@38874.8]
  wire  _T_93359; // @[LoadQueue.scala 233:86:@38875.8]
  wire  _T_93360; // @[LoadQueue.scala 233:86:@38876.8]
  wire  _T_93361; // @[LoadQueue.scala 233:86:@38877.8]
  wire  _T_93362; // @[LoadQueue.scala 233:86:@38878.8]
  wire  _T_93363; // @[LoadQueue.scala 233:86:@38879.8]
  wire  _T_93364; // @[LoadQueue.scala 233:86:@38880.8]
  wire  _T_93365; // @[LoadQueue.scala 233:86:@38881.8]
  wire  _T_93366; // @[LoadQueue.scala 233:86:@38882.8]
  wire  _T_93367; // @[LoadQueue.scala 233:86:@38883.8]
  wire  _T_93368; // @[LoadQueue.scala 233:86:@38884.8]
  wire  _T_93369; // @[LoadQueue.scala 233:86:@38885.8]
  wire  _T_93370; // @[LoadQueue.scala 233:86:@38886.8]
  wire  _T_93372; // @[LoadQueue.scala 233:38:@38887.8]
  wire  _T_93391; // @[LoadQueue.scala 234:11:@38904.8]
  wire  _T_93392; // @[LoadQueue.scala 233:103:@38905.8]
  wire  _GEN_2020; // @[LoadQueue.scala 230:110:@38870.6]
  wire  loadRequest_13; // @[LoadQueue.scala 229:71:@38864.4]
  wire [15:0] _T_90458; // @[Mux.scala 31:69:@36523.4]
  wire  _T_93260; // @[LoadQueue.scala 229:41:@38780.4]
  wire  _T_93261; // @[LoadQueue.scala 229:38:@38781.4]
  wire  _T_93263; // @[LoadQueue.scala 230:12:@38783.6]
  reg  prevPriorityRequest_12; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_742;
  wire  _T_93265; // @[LoadQueue.scala 230:46:@38784.6]
  wire  _T_93266; // @[LoadQueue.scala 230:43:@38785.6]
  wire  _T_93268; // @[LoadQueue.scala 230:84:@38786.6]
  wire  _T_93269; // @[LoadQueue.scala 230:81:@38787.6]
  wire  _T_93272; // @[LoadQueue.scala 233:86:@38790.8]
  wire  _T_93273; // @[LoadQueue.scala 233:86:@38791.8]
  wire  _T_93274; // @[LoadQueue.scala 233:86:@38792.8]
  wire  _T_93275; // @[LoadQueue.scala 233:86:@38793.8]
  wire  _T_93276; // @[LoadQueue.scala 233:86:@38794.8]
  wire  _T_93277; // @[LoadQueue.scala 233:86:@38795.8]
  wire  _T_93278; // @[LoadQueue.scala 233:86:@38796.8]
  wire  _T_93279; // @[LoadQueue.scala 233:86:@38797.8]
  wire  _T_93280; // @[LoadQueue.scala 233:86:@38798.8]
  wire  _T_93281; // @[LoadQueue.scala 233:86:@38799.8]
  wire  _T_93282; // @[LoadQueue.scala 233:86:@38800.8]
  wire  _T_93283; // @[LoadQueue.scala 233:86:@38801.8]
  wire  _T_93284; // @[LoadQueue.scala 233:86:@38802.8]
  wire  _T_93285; // @[LoadQueue.scala 233:86:@38803.8]
  wire  _T_93286; // @[LoadQueue.scala 233:86:@38804.8]
  wire  _T_93288; // @[LoadQueue.scala 233:38:@38805.8]
  wire  _T_93307; // @[LoadQueue.scala 234:11:@38822.8]
  wire  _T_93308; // @[LoadQueue.scala 233:103:@38823.8]
  wire  _GEN_2016; // @[LoadQueue.scala 230:110:@38788.6]
  wire  loadRequest_12; // @[LoadQueue.scala 229:71:@38782.4]
  wire [15:0] _T_90459; // @[Mux.scala 31:69:@36524.4]
  wire  _T_93176; // @[LoadQueue.scala 229:41:@38698.4]
  wire  _T_93177; // @[LoadQueue.scala 229:38:@38699.4]
  wire  _T_93179; // @[LoadQueue.scala 230:12:@38701.6]
  reg  prevPriorityRequest_11; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_743;
  wire  _T_93181; // @[LoadQueue.scala 230:46:@38702.6]
  wire  _T_93182; // @[LoadQueue.scala 230:43:@38703.6]
  wire  _T_93184; // @[LoadQueue.scala 230:84:@38704.6]
  wire  _T_93185; // @[LoadQueue.scala 230:81:@38705.6]
  wire  _T_93188; // @[LoadQueue.scala 233:86:@38708.8]
  wire  _T_93189; // @[LoadQueue.scala 233:86:@38709.8]
  wire  _T_93190; // @[LoadQueue.scala 233:86:@38710.8]
  wire  _T_93191; // @[LoadQueue.scala 233:86:@38711.8]
  wire  _T_93192; // @[LoadQueue.scala 233:86:@38712.8]
  wire  _T_93193; // @[LoadQueue.scala 233:86:@38713.8]
  wire  _T_93194; // @[LoadQueue.scala 233:86:@38714.8]
  wire  _T_93195; // @[LoadQueue.scala 233:86:@38715.8]
  wire  _T_93196; // @[LoadQueue.scala 233:86:@38716.8]
  wire  _T_93197; // @[LoadQueue.scala 233:86:@38717.8]
  wire  _T_93198; // @[LoadQueue.scala 233:86:@38718.8]
  wire  _T_93199; // @[LoadQueue.scala 233:86:@38719.8]
  wire  _T_93200; // @[LoadQueue.scala 233:86:@38720.8]
  wire  _T_93201; // @[LoadQueue.scala 233:86:@38721.8]
  wire  _T_93202; // @[LoadQueue.scala 233:86:@38722.8]
  wire  _T_93204; // @[LoadQueue.scala 233:38:@38723.8]
  wire  _T_93223; // @[LoadQueue.scala 234:11:@38740.8]
  wire  _T_93224; // @[LoadQueue.scala 233:103:@38741.8]
  wire  _GEN_2012; // @[LoadQueue.scala 230:110:@38706.6]
  wire  loadRequest_11; // @[LoadQueue.scala 229:71:@38700.4]
  wire [15:0] _T_90460; // @[Mux.scala 31:69:@36525.4]
  wire  _T_93092; // @[LoadQueue.scala 229:41:@38616.4]
  wire  _T_93093; // @[LoadQueue.scala 229:38:@38617.4]
  wire  _T_93095; // @[LoadQueue.scala 230:12:@38619.6]
  reg  prevPriorityRequest_10; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_744;
  wire  _T_93097; // @[LoadQueue.scala 230:46:@38620.6]
  wire  _T_93098; // @[LoadQueue.scala 230:43:@38621.6]
  wire  _T_93100; // @[LoadQueue.scala 230:84:@38622.6]
  wire  _T_93101; // @[LoadQueue.scala 230:81:@38623.6]
  wire  _T_93104; // @[LoadQueue.scala 233:86:@38626.8]
  wire  _T_93105; // @[LoadQueue.scala 233:86:@38627.8]
  wire  _T_93106; // @[LoadQueue.scala 233:86:@38628.8]
  wire  _T_93107; // @[LoadQueue.scala 233:86:@38629.8]
  wire  _T_93108; // @[LoadQueue.scala 233:86:@38630.8]
  wire  _T_93109; // @[LoadQueue.scala 233:86:@38631.8]
  wire  _T_93110; // @[LoadQueue.scala 233:86:@38632.8]
  wire  _T_93111; // @[LoadQueue.scala 233:86:@38633.8]
  wire  _T_93112; // @[LoadQueue.scala 233:86:@38634.8]
  wire  _T_93113; // @[LoadQueue.scala 233:86:@38635.8]
  wire  _T_93114; // @[LoadQueue.scala 233:86:@38636.8]
  wire  _T_93115; // @[LoadQueue.scala 233:86:@38637.8]
  wire  _T_93116; // @[LoadQueue.scala 233:86:@38638.8]
  wire  _T_93117; // @[LoadQueue.scala 233:86:@38639.8]
  wire  _T_93118; // @[LoadQueue.scala 233:86:@38640.8]
  wire  _T_93120; // @[LoadQueue.scala 233:38:@38641.8]
  wire  _T_93139; // @[LoadQueue.scala 234:11:@38658.8]
  wire  _T_93140; // @[LoadQueue.scala 233:103:@38659.8]
  wire  _GEN_2008; // @[LoadQueue.scala 230:110:@38624.6]
  wire  loadRequest_10; // @[LoadQueue.scala 229:71:@38618.4]
  wire [15:0] _T_90461; // @[Mux.scala 31:69:@36526.4]
  wire  _T_93008; // @[LoadQueue.scala 229:41:@38534.4]
  wire  _T_93009; // @[LoadQueue.scala 229:38:@38535.4]
  wire  _T_93011; // @[LoadQueue.scala 230:12:@38537.6]
  reg  prevPriorityRequest_9; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_745;
  wire  _T_93013; // @[LoadQueue.scala 230:46:@38538.6]
  wire  _T_93014; // @[LoadQueue.scala 230:43:@38539.6]
  wire  _T_93016; // @[LoadQueue.scala 230:84:@38540.6]
  wire  _T_93017; // @[LoadQueue.scala 230:81:@38541.6]
  wire  _T_93020; // @[LoadQueue.scala 233:86:@38544.8]
  wire  _T_93021; // @[LoadQueue.scala 233:86:@38545.8]
  wire  _T_93022; // @[LoadQueue.scala 233:86:@38546.8]
  wire  _T_93023; // @[LoadQueue.scala 233:86:@38547.8]
  wire  _T_93024; // @[LoadQueue.scala 233:86:@38548.8]
  wire  _T_93025; // @[LoadQueue.scala 233:86:@38549.8]
  wire  _T_93026; // @[LoadQueue.scala 233:86:@38550.8]
  wire  _T_93027; // @[LoadQueue.scala 233:86:@38551.8]
  wire  _T_93028; // @[LoadQueue.scala 233:86:@38552.8]
  wire  _T_93029; // @[LoadQueue.scala 233:86:@38553.8]
  wire  _T_93030; // @[LoadQueue.scala 233:86:@38554.8]
  wire  _T_93031; // @[LoadQueue.scala 233:86:@38555.8]
  wire  _T_93032; // @[LoadQueue.scala 233:86:@38556.8]
  wire  _T_93033; // @[LoadQueue.scala 233:86:@38557.8]
  wire  _T_93034; // @[LoadQueue.scala 233:86:@38558.8]
  wire  _T_93036; // @[LoadQueue.scala 233:38:@38559.8]
  wire  _T_93055; // @[LoadQueue.scala 234:11:@38576.8]
  wire  _T_93056; // @[LoadQueue.scala 233:103:@38577.8]
  wire  _GEN_2004; // @[LoadQueue.scala 230:110:@38542.6]
  wire  loadRequest_9; // @[LoadQueue.scala 229:71:@38536.4]
  wire [15:0] _T_90462; // @[Mux.scala 31:69:@36527.4]
  wire  _T_92924; // @[LoadQueue.scala 229:41:@38452.4]
  wire  _T_92925; // @[LoadQueue.scala 229:38:@38453.4]
  wire  _T_92927; // @[LoadQueue.scala 230:12:@38455.6]
  reg  prevPriorityRequest_8; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_746;
  wire  _T_92929; // @[LoadQueue.scala 230:46:@38456.6]
  wire  _T_92930; // @[LoadQueue.scala 230:43:@38457.6]
  wire  _T_92932; // @[LoadQueue.scala 230:84:@38458.6]
  wire  _T_92933; // @[LoadQueue.scala 230:81:@38459.6]
  wire  _T_92936; // @[LoadQueue.scala 233:86:@38462.8]
  wire  _T_92937; // @[LoadQueue.scala 233:86:@38463.8]
  wire  _T_92938; // @[LoadQueue.scala 233:86:@38464.8]
  wire  _T_92939; // @[LoadQueue.scala 233:86:@38465.8]
  wire  _T_92940; // @[LoadQueue.scala 233:86:@38466.8]
  wire  _T_92941; // @[LoadQueue.scala 233:86:@38467.8]
  wire  _T_92942; // @[LoadQueue.scala 233:86:@38468.8]
  wire  _T_92943; // @[LoadQueue.scala 233:86:@38469.8]
  wire  _T_92944; // @[LoadQueue.scala 233:86:@38470.8]
  wire  _T_92945; // @[LoadQueue.scala 233:86:@38471.8]
  wire  _T_92946; // @[LoadQueue.scala 233:86:@38472.8]
  wire  _T_92947; // @[LoadQueue.scala 233:86:@38473.8]
  wire  _T_92948; // @[LoadQueue.scala 233:86:@38474.8]
  wire  _T_92949; // @[LoadQueue.scala 233:86:@38475.8]
  wire  _T_92950; // @[LoadQueue.scala 233:86:@38476.8]
  wire  _T_92952; // @[LoadQueue.scala 233:38:@38477.8]
  wire  _T_92971; // @[LoadQueue.scala 234:11:@38494.8]
  wire  _T_92972; // @[LoadQueue.scala 233:103:@38495.8]
  wire  _GEN_2000; // @[LoadQueue.scala 230:110:@38460.6]
  wire  loadRequest_8; // @[LoadQueue.scala 229:71:@38454.4]
  wire [15:0] _T_90463; // @[Mux.scala 31:69:@36528.4]
  wire  _T_92840; // @[LoadQueue.scala 229:41:@38370.4]
  wire  _T_92841; // @[LoadQueue.scala 229:38:@38371.4]
  wire  _T_92843; // @[LoadQueue.scala 230:12:@38373.6]
  reg  prevPriorityRequest_7; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_747;
  wire  _T_92845; // @[LoadQueue.scala 230:46:@38374.6]
  wire  _T_92846; // @[LoadQueue.scala 230:43:@38375.6]
  wire  _T_92848; // @[LoadQueue.scala 230:84:@38376.6]
  wire  _T_92849; // @[LoadQueue.scala 230:81:@38377.6]
  wire  _T_92852; // @[LoadQueue.scala 233:86:@38380.8]
  wire  _T_92853; // @[LoadQueue.scala 233:86:@38381.8]
  wire  _T_92854; // @[LoadQueue.scala 233:86:@38382.8]
  wire  _T_92855; // @[LoadQueue.scala 233:86:@38383.8]
  wire  _T_92856; // @[LoadQueue.scala 233:86:@38384.8]
  wire  _T_92857; // @[LoadQueue.scala 233:86:@38385.8]
  wire  _T_92858; // @[LoadQueue.scala 233:86:@38386.8]
  wire  _T_92859; // @[LoadQueue.scala 233:86:@38387.8]
  wire  _T_92860; // @[LoadQueue.scala 233:86:@38388.8]
  wire  _T_92861; // @[LoadQueue.scala 233:86:@38389.8]
  wire  _T_92862; // @[LoadQueue.scala 233:86:@38390.8]
  wire  _T_92863; // @[LoadQueue.scala 233:86:@38391.8]
  wire  _T_92864; // @[LoadQueue.scala 233:86:@38392.8]
  wire  _T_92865; // @[LoadQueue.scala 233:86:@38393.8]
  wire  _T_92866; // @[LoadQueue.scala 233:86:@38394.8]
  wire  _T_92868; // @[LoadQueue.scala 233:38:@38395.8]
  wire  _T_92887; // @[LoadQueue.scala 234:11:@38412.8]
  wire  _T_92888; // @[LoadQueue.scala 233:103:@38413.8]
  wire  _GEN_1996; // @[LoadQueue.scala 230:110:@38378.6]
  wire  loadRequest_7; // @[LoadQueue.scala 229:71:@38372.4]
  wire [15:0] _T_90464; // @[Mux.scala 31:69:@36529.4]
  wire  _T_92756; // @[LoadQueue.scala 229:41:@38288.4]
  wire  _T_92757; // @[LoadQueue.scala 229:38:@38289.4]
  wire  _T_92759; // @[LoadQueue.scala 230:12:@38291.6]
  reg  prevPriorityRequest_6; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_748;
  wire  _T_92761; // @[LoadQueue.scala 230:46:@38292.6]
  wire  _T_92762; // @[LoadQueue.scala 230:43:@38293.6]
  wire  _T_92764; // @[LoadQueue.scala 230:84:@38294.6]
  wire  _T_92765; // @[LoadQueue.scala 230:81:@38295.6]
  wire  _T_92768; // @[LoadQueue.scala 233:86:@38298.8]
  wire  _T_92769; // @[LoadQueue.scala 233:86:@38299.8]
  wire  _T_92770; // @[LoadQueue.scala 233:86:@38300.8]
  wire  _T_92771; // @[LoadQueue.scala 233:86:@38301.8]
  wire  _T_92772; // @[LoadQueue.scala 233:86:@38302.8]
  wire  _T_92773; // @[LoadQueue.scala 233:86:@38303.8]
  wire  _T_92774; // @[LoadQueue.scala 233:86:@38304.8]
  wire  _T_92775; // @[LoadQueue.scala 233:86:@38305.8]
  wire  _T_92776; // @[LoadQueue.scala 233:86:@38306.8]
  wire  _T_92777; // @[LoadQueue.scala 233:86:@38307.8]
  wire  _T_92778; // @[LoadQueue.scala 233:86:@38308.8]
  wire  _T_92779; // @[LoadQueue.scala 233:86:@38309.8]
  wire  _T_92780; // @[LoadQueue.scala 233:86:@38310.8]
  wire  _T_92781; // @[LoadQueue.scala 233:86:@38311.8]
  wire  _T_92782; // @[LoadQueue.scala 233:86:@38312.8]
  wire  _T_92784; // @[LoadQueue.scala 233:38:@38313.8]
  wire  _T_92803; // @[LoadQueue.scala 234:11:@38330.8]
  wire  _T_92804; // @[LoadQueue.scala 233:103:@38331.8]
  wire  _GEN_1992; // @[LoadQueue.scala 230:110:@38296.6]
  wire  loadRequest_6; // @[LoadQueue.scala 229:71:@38290.4]
  wire [15:0] _T_90465; // @[Mux.scala 31:69:@36530.4]
  wire  _T_92672; // @[LoadQueue.scala 229:41:@38206.4]
  wire  _T_92673; // @[LoadQueue.scala 229:38:@38207.4]
  wire  _T_92675; // @[LoadQueue.scala 230:12:@38209.6]
  reg  prevPriorityRequest_5; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_749;
  wire  _T_92677; // @[LoadQueue.scala 230:46:@38210.6]
  wire  _T_92678; // @[LoadQueue.scala 230:43:@38211.6]
  wire  _T_92680; // @[LoadQueue.scala 230:84:@38212.6]
  wire  _T_92681; // @[LoadQueue.scala 230:81:@38213.6]
  wire  _T_92684; // @[LoadQueue.scala 233:86:@38216.8]
  wire  _T_92685; // @[LoadQueue.scala 233:86:@38217.8]
  wire  _T_92686; // @[LoadQueue.scala 233:86:@38218.8]
  wire  _T_92687; // @[LoadQueue.scala 233:86:@38219.8]
  wire  _T_92688; // @[LoadQueue.scala 233:86:@38220.8]
  wire  _T_92689; // @[LoadQueue.scala 233:86:@38221.8]
  wire  _T_92690; // @[LoadQueue.scala 233:86:@38222.8]
  wire  _T_92691; // @[LoadQueue.scala 233:86:@38223.8]
  wire  _T_92692; // @[LoadQueue.scala 233:86:@38224.8]
  wire  _T_92693; // @[LoadQueue.scala 233:86:@38225.8]
  wire  _T_92694; // @[LoadQueue.scala 233:86:@38226.8]
  wire  _T_92695; // @[LoadQueue.scala 233:86:@38227.8]
  wire  _T_92696; // @[LoadQueue.scala 233:86:@38228.8]
  wire  _T_92697; // @[LoadQueue.scala 233:86:@38229.8]
  wire  _T_92698; // @[LoadQueue.scala 233:86:@38230.8]
  wire  _T_92700; // @[LoadQueue.scala 233:38:@38231.8]
  wire  _T_92719; // @[LoadQueue.scala 234:11:@38248.8]
  wire  _T_92720; // @[LoadQueue.scala 233:103:@38249.8]
  wire  _GEN_1988; // @[LoadQueue.scala 230:110:@38214.6]
  wire  loadRequest_5; // @[LoadQueue.scala 229:71:@38208.4]
  wire [15:0] _T_90466; // @[Mux.scala 31:69:@36531.4]
  wire  _T_92588; // @[LoadQueue.scala 229:41:@38124.4]
  wire  _T_92589; // @[LoadQueue.scala 229:38:@38125.4]
  wire  _T_92591; // @[LoadQueue.scala 230:12:@38127.6]
  reg  prevPriorityRequest_4; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_750;
  wire  _T_92593; // @[LoadQueue.scala 230:46:@38128.6]
  wire  _T_92594; // @[LoadQueue.scala 230:43:@38129.6]
  wire  _T_92596; // @[LoadQueue.scala 230:84:@38130.6]
  wire  _T_92597; // @[LoadQueue.scala 230:81:@38131.6]
  wire  _T_92600; // @[LoadQueue.scala 233:86:@38134.8]
  wire  _T_92601; // @[LoadQueue.scala 233:86:@38135.8]
  wire  _T_92602; // @[LoadQueue.scala 233:86:@38136.8]
  wire  _T_92603; // @[LoadQueue.scala 233:86:@38137.8]
  wire  _T_92604; // @[LoadQueue.scala 233:86:@38138.8]
  wire  _T_92605; // @[LoadQueue.scala 233:86:@38139.8]
  wire  _T_92606; // @[LoadQueue.scala 233:86:@38140.8]
  wire  _T_92607; // @[LoadQueue.scala 233:86:@38141.8]
  wire  _T_92608; // @[LoadQueue.scala 233:86:@38142.8]
  wire  _T_92609; // @[LoadQueue.scala 233:86:@38143.8]
  wire  _T_92610; // @[LoadQueue.scala 233:86:@38144.8]
  wire  _T_92611; // @[LoadQueue.scala 233:86:@38145.8]
  wire  _T_92612; // @[LoadQueue.scala 233:86:@38146.8]
  wire  _T_92613; // @[LoadQueue.scala 233:86:@38147.8]
  wire  _T_92614; // @[LoadQueue.scala 233:86:@38148.8]
  wire  _T_92616; // @[LoadQueue.scala 233:38:@38149.8]
  wire  _T_92635; // @[LoadQueue.scala 234:11:@38166.8]
  wire  _T_92636; // @[LoadQueue.scala 233:103:@38167.8]
  wire  _GEN_1984; // @[LoadQueue.scala 230:110:@38132.6]
  wire  loadRequest_4; // @[LoadQueue.scala 229:71:@38126.4]
  wire [15:0] _T_90467; // @[Mux.scala 31:69:@36532.4]
  wire  _T_92504; // @[LoadQueue.scala 229:41:@38042.4]
  wire  _T_92505; // @[LoadQueue.scala 229:38:@38043.4]
  wire  _T_92507; // @[LoadQueue.scala 230:12:@38045.6]
  reg  prevPriorityRequest_3; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_751;
  wire  _T_92509; // @[LoadQueue.scala 230:46:@38046.6]
  wire  _T_92510; // @[LoadQueue.scala 230:43:@38047.6]
  wire  _T_92512; // @[LoadQueue.scala 230:84:@38048.6]
  wire  _T_92513; // @[LoadQueue.scala 230:81:@38049.6]
  wire  _T_92516; // @[LoadQueue.scala 233:86:@38052.8]
  wire  _T_92517; // @[LoadQueue.scala 233:86:@38053.8]
  wire  _T_92518; // @[LoadQueue.scala 233:86:@38054.8]
  wire  _T_92519; // @[LoadQueue.scala 233:86:@38055.8]
  wire  _T_92520; // @[LoadQueue.scala 233:86:@38056.8]
  wire  _T_92521; // @[LoadQueue.scala 233:86:@38057.8]
  wire  _T_92522; // @[LoadQueue.scala 233:86:@38058.8]
  wire  _T_92523; // @[LoadQueue.scala 233:86:@38059.8]
  wire  _T_92524; // @[LoadQueue.scala 233:86:@38060.8]
  wire  _T_92525; // @[LoadQueue.scala 233:86:@38061.8]
  wire  _T_92526; // @[LoadQueue.scala 233:86:@38062.8]
  wire  _T_92527; // @[LoadQueue.scala 233:86:@38063.8]
  wire  _T_92528; // @[LoadQueue.scala 233:86:@38064.8]
  wire  _T_92529; // @[LoadQueue.scala 233:86:@38065.8]
  wire  _T_92530; // @[LoadQueue.scala 233:86:@38066.8]
  wire  _T_92532; // @[LoadQueue.scala 233:38:@38067.8]
  wire  _T_92551; // @[LoadQueue.scala 234:11:@38084.8]
  wire  _T_92552; // @[LoadQueue.scala 233:103:@38085.8]
  wire  _GEN_1980; // @[LoadQueue.scala 230:110:@38050.6]
  wire  loadRequest_3; // @[LoadQueue.scala 229:71:@38044.4]
  wire [15:0] _T_90468; // @[Mux.scala 31:69:@36533.4]
  wire  _T_92420; // @[LoadQueue.scala 229:41:@37960.4]
  wire  _T_92421; // @[LoadQueue.scala 229:38:@37961.4]
  wire  _T_92423; // @[LoadQueue.scala 230:12:@37963.6]
  reg  prevPriorityRequest_2; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_752;
  wire  _T_92425; // @[LoadQueue.scala 230:46:@37964.6]
  wire  _T_92426; // @[LoadQueue.scala 230:43:@37965.6]
  wire  _T_92428; // @[LoadQueue.scala 230:84:@37966.6]
  wire  _T_92429; // @[LoadQueue.scala 230:81:@37967.6]
  wire  _T_92432; // @[LoadQueue.scala 233:86:@37970.8]
  wire  _T_92433; // @[LoadQueue.scala 233:86:@37971.8]
  wire  _T_92434; // @[LoadQueue.scala 233:86:@37972.8]
  wire  _T_92435; // @[LoadQueue.scala 233:86:@37973.8]
  wire  _T_92436; // @[LoadQueue.scala 233:86:@37974.8]
  wire  _T_92437; // @[LoadQueue.scala 233:86:@37975.8]
  wire  _T_92438; // @[LoadQueue.scala 233:86:@37976.8]
  wire  _T_92439; // @[LoadQueue.scala 233:86:@37977.8]
  wire  _T_92440; // @[LoadQueue.scala 233:86:@37978.8]
  wire  _T_92441; // @[LoadQueue.scala 233:86:@37979.8]
  wire  _T_92442; // @[LoadQueue.scala 233:86:@37980.8]
  wire  _T_92443; // @[LoadQueue.scala 233:86:@37981.8]
  wire  _T_92444; // @[LoadQueue.scala 233:86:@37982.8]
  wire  _T_92445; // @[LoadQueue.scala 233:86:@37983.8]
  wire  _T_92446; // @[LoadQueue.scala 233:86:@37984.8]
  wire  _T_92448; // @[LoadQueue.scala 233:38:@37985.8]
  wire  _T_92467; // @[LoadQueue.scala 234:11:@38002.8]
  wire  _T_92468; // @[LoadQueue.scala 233:103:@38003.8]
  wire  _GEN_1976; // @[LoadQueue.scala 230:110:@37968.6]
  wire  loadRequest_2; // @[LoadQueue.scala 229:71:@37962.4]
  wire [15:0] _T_90469; // @[Mux.scala 31:69:@36534.4]
  wire  _T_92336; // @[LoadQueue.scala 229:41:@37878.4]
  wire  _T_92337; // @[LoadQueue.scala 229:38:@37879.4]
  wire  _T_92339; // @[LoadQueue.scala 230:12:@37881.6]
  reg  prevPriorityRequest_1; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_753;
  wire  _T_92341; // @[LoadQueue.scala 230:46:@37882.6]
  wire  _T_92342; // @[LoadQueue.scala 230:43:@37883.6]
  wire  _T_92344; // @[LoadQueue.scala 230:84:@37884.6]
  wire  _T_92345; // @[LoadQueue.scala 230:81:@37885.6]
  wire  _T_92348; // @[LoadQueue.scala 233:86:@37888.8]
  wire  _T_92349; // @[LoadQueue.scala 233:86:@37889.8]
  wire  _T_92350; // @[LoadQueue.scala 233:86:@37890.8]
  wire  _T_92351; // @[LoadQueue.scala 233:86:@37891.8]
  wire  _T_92352; // @[LoadQueue.scala 233:86:@37892.8]
  wire  _T_92353; // @[LoadQueue.scala 233:86:@37893.8]
  wire  _T_92354; // @[LoadQueue.scala 233:86:@37894.8]
  wire  _T_92355; // @[LoadQueue.scala 233:86:@37895.8]
  wire  _T_92356; // @[LoadQueue.scala 233:86:@37896.8]
  wire  _T_92357; // @[LoadQueue.scala 233:86:@37897.8]
  wire  _T_92358; // @[LoadQueue.scala 233:86:@37898.8]
  wire  _T_92359; // @[LoadQueue.scala 233:86:@37899.8]
  wire  _T_92360; // @[LoadQueue.scala 233:86:@37900.8]
  wire  _T_92361; // @[LoadQueue.scala 233:86:@37901.8]
  wire  _T_92362; // @[LoadQueue.scala 233:86:@37902.8]
  wire  _T_92364; // @[LoadQueue.scala 233:38:@37903.8]
  wire  _T_92383; // @[LoadQueue.scala 234:11:@37920.8]
  wire  _T_92384; // @[LoadQueue.scala 233:103:@37921.8]
  wire  _GEN_1972; // @[LoadQueue.scala 230:110:@37886.6]
  wire  loadRequest_1; // @[LoadQueue.scala 229:71:@37880.4]
  wire [15:0] _T_90470; // @[Mux.scala 31:69:@36535.4]
  wire  _T_92252; // @[LoadQueue.scala 229:41:@37796.4]
  wire  _T_92253; // @[LoadQueue.scala 229:38:@37797.4]
  wire  _T_92255; // @[LoadQueue.scala 230:12:@37799.6]
  reg  prevPriorityRequest_0; // @[LoadQueue.scala 207:36:@37628.4]
  reg [31:0] _RAND_754;
  wire  _T_92257; // @[LoadQueue.scala 230:46:@37800.6]
  wire  _T_92258; // @[LoadQueue.scala 230:43:@37801.6]
  wire  _T_92260; // @[LoadQueue.scala 230:84:@37802.6]
  wire  _T_92261; // @[LoadQueue.scala 230:81:@37803.6]
  wire  _T_92264; // @[LoadQueue.scala 233:86:@37806.8]
  wire  _T_92265; // @[LoadQueue.scala 233:86:@37807.8]
  wire  _T_92266; // @[LoadQueue.scala 233:86:@37808.8]
  wire  _T_92267; // @[LoadQueue.scala 233:86:@37809.8]
  wire  _T_92268; // @[LoadQueue.scala 233:86:@37810.8]
  wire  _T_92269; // @[LoadQueue.scala 233:86:@37811.8]
  wire  _T_92270; // @[LoadQueue.scala 233:86:@37812.8]
  wire  _T_92271; // @[LoadQueue.scala 233:86:@37813.8]
  wire  _T_92272; // @[LoadQueue.scala 233:86:@37814.8]
  wire  _T_92273; // @[LoadQueue.scala 233:86:@37815.8]
  wire  _T_92274; // @[LoadQueue.scala 233:86:@37816.8]
  wire  _T_92275; // @[LoadQueue.scala 233:86:@37817.8]
  wire  _T_92276; // @[LoadQueue.scala 233:86:@37818.8]
  wire  _T_92277; // @[LoadQueue.scala 233:86:@37819.8]
  wire  _T_92278; // @[LoadQueue.scala 233:86:@37820.8]
  wire  _T_92280; // @[LoadQueue.scala 233:38:@37821.8]
  wire  _T_92299; // @[LoadQueue.scala 234:11:@37838.8]
  wire  _T_92300; // @[LoadQueue.scala 233:103:@37839.8]
  wire  _GEN_1968; // @[LoadQueue.scala 230:110:@37804.6]
  wire  loadRequest_0; // @[LoadQueue.scala 229:71:@37798.4]
  wire [15:0] _T_90471; // @[Mux.scala 31:69:@36536.4]
  wire  _T_90472; // @[OneHot.scala 66:30:@36537.4]
  wire  _T_90473; // @[OneHot.scala 66:30:@36538.4]
  wire  _T_90474; // @[OneHot.scala 66:30:@36539.4]
  wire  _T_90475; // @[OneHot.scala 66:30:@36540.4]
  wire  _T_90476; // @[OneHot.scala 66:30:@36541.4]
  wire  _T_90477; // @[OneHot.scala 66:30:@36542.4]
  wire  _T_90478; // @[OneHot.scala 66:30:@36543.4]
  wire  _T_90479; // @[OneHot.scala 66:30:@36544.4]
  wire  _T_90480; // @[OneHot.scala 66:30:@36545.4]
  wire  _T_90481; // @[OneHot.scala 66:30:@36546.4]
  wire  _T_90482; // @[OneHot.scala 66:30:@36547.4]
  wire  _T_90483; // @[OneHot.scala 66:30:@36548.4]
  wire  _T_90484; // @[OneHot.scala 66:30:@36549.4]
  wire  _T_90485; // @[OneHot.scala 66:30:@36550.4]
  wire  _T_90486; // @[OneHot.scala 66:30:@36551.4]
  wire  _T_90487; // @[OneHot.scala 66:30:@36552.4]
  wire [15:0] _T_90528; // @[Mux.scala 31:69:@36570.4]
  wire [15:0] _T_90529; // @[Mux.scala 31:69:@36571.4]
  wire [15:0] _T_90530; // @[Mux.scala 31:69:@36572.4]
  wire [15:0] _T_90531; // @[Mux.scala 31:69:@36573.4]
  wire [15:0] _T_90532; // @[Mux.scala 31:69:@36574.4]
  wire [15:0] _T_90533; // @[Mux.scala 31:69:@36575.4]
  wire [15:0] _T_90534; // @[Mux.scala 31:69:@36576.4]
  wire [15:0] _T_90535; // @[Mux.scala 31:69:@36577.4]
  wire [15:0] _T_90536; // @[Mux.scala 31:69:@36578.4]
  wire [15:0] _T_90537; // @[Mux.scala 31:69:@36579.4]
  wire [15:0] _T_90538; // @[Mux.scala 31:69:@36580.4]
  wire [15:0] _T_90539; // @[Mux.scala 31:69:@36581.4]
  wire [15:0] _T_90540; // @[Mux.scala 31:69:@36582.4]
  wire [15:0] _T_90541; // @[Mux.scala 31:69:@36583.4]
  wire [15:0] _T_90542; // @[Mux.scala 31:69:@36584.4]
  wire [15:0] _T_90543; // @[Mux.scala 31:69:@36585.4]
  wire  _T_90544; // @[OneHot.scala 66:30:@36586.4]
  wire  _T_90545; // @[OneHot.scala 66:30:@36587.4]
  wire  _T_90546; // @[OneHot.scala 66:30:@36588.4]
  wire  _T_90547; // @[OneHot.scala 66:30:@36589.4]
  wire  _T_90548; // @[OneHot.scala 66:30:@36590.4]
  wire  _T_90549; // @[OneHot.scala 66:30:@36591.4]
  wire  _T_90550; // @[OneHot.scala 66:30:@36592.4]
  wire  _T_90551; // @[OneHot.scala 66:30:@36593.4]
  wire  _T_90552; // @[OneHot.scala 66:30:@36594.4]
  wire  _T_90553; // @[OneHot.scala 66:30:@36595.4]
  wire  _T_90554; // @[OneHot.scala 66:30:@36596.4]
  wire  _T_90555; // @[OneHot.scala 66:30:@36597.4]
  wire  _T_90556; // @[OneHot.scala 66:30:@36598.4]
  wire  _T_90557; // @[OneHot.scala 66:30:@36599.4]
  wire  _T_90558; // @[OneHot.scala 66:30:@36600.4]
  wire  _T_90559; // @[OneHot.scala 66:30:@36601.4]
  wire [15:0] _T_90600; // @[Mux.scala 31:69:@36619.4]
  wire [15:0] _T_90601; // @[Mux.scala 31:69:@36620.4]
  wire [15:0] _T_90602; // @[Mux.scala 31:69:@36621.4]
  wire [15:0] _T_90603; // @[Mux.scala 31:69:@36622.4]
  wire [15:0] _T_90604; // @[Mux.scala 31:69:@36623.4]
  wire [15:0] _T_90605; // @[Mux.scala 31:69:@36624.4]
  wire [15:0] _T_90606; // @[Mux.scala 31:69:@36625.4]
  wire [15:0] _T_90607; // @[Mux.scala 31:69:@36626.4]
  wire [15:0] _T_90608; // @[Mux.scala 31:69:@36627.4]
  wire [15:0] _T_90609; // @[Mux.scala 31:69:@36628.4]
  wire [15:0] _T_90610; // @[Mux.scala 31:69:@36629.4]
  wire [15:0] _T_90611; // @[Mux.scala 31:69:@36630.4]
  wire [15:0] _T_90612; // @[Mux.scala 31:69:@36631.4]
  wire [15:0] _T_90613; // @[Mux.scala 31:69:@36632.4]
  wire [15:0] _T_90614; // @[Mux.scala 31:69:@36633.4]
  wire [15:0] _T_90615; // @[Mux.scala 31:69:@36634.4]
  wire  _T_90616; // @[OneHot.scala 66:30:@36635.4]
  wire  _T_90617; // @[OneHot.scala 66:30:@36636.4]
  wire  _T_90618; // @[OneHot.scala 66:30:@36637.4]
  wire  _T_90619; // @[OneHot.scala 66:30:@36638.4]
  wire  _T_90620; // @[OneHot.scala 66:30:@36639.4]
  wire  _T_90621; // @[OneHot.scala 66:30:@36640.4]
  wire  _T_90622; // @[OneHot.scala 66:30:@36641.4]
  wire  _T_90623; // @[OneHot.scala 66:30:@36642.4]
  wire  _T_90624; // @[OneHot.scala 66:30:@36643.4]
  wire  _T_90625; // @[OneHot.scala 66:30:@36644.4]
  wire  _T_90626; // @[OneHot.scala 66:30:@36645.4]
  wire  _T_90627; // @[OneHot.scala 66:30:@36646.4]
  wire  _T_90628; // @[OneHot.scala 66:30:@36647.4]
  wire  _T_90629; // @[OneHot.scala 66:30:@36648.4]
  wire  _T_90630; // @[OneHot.scala 66:30:@36649.4]
  wire  _T_90631; // @[OneHot.scala 66:30:@36650.4]
  wire [15:0] _T_90672; // @[Mux.scala 31:69:@36668.4]
  wire [15:0] _T_90673; // @[Mux.scala 31:69:@36669.4]
  wire [15:0] _T_90674; // @[Mux.scala 31:69:@36670.4]
  wire [15:0] _T_90675; // @[Mux.scala 31:69:@36671.4]
  wire [15:0] _T_90676; // @[Mux.scala 31:69:@36672.4]
  wire [15:0] _T_90677; // @[Mux.scala 31:69:@36673.4]
  wire [15:0] _T_90678; // @[Mux.scala 31:69:@36674.4]
  wire [15:0] _T_90679; // @[Mux.scala 31:69:@36675.4]
  wire [15:0] _T_90680; // @[Mux.scala 31:69:@36676.4]
  wire [15:0] _T_90681; // @[Mux.scala 31:69:@36677.4]
  wire [15:0] _T_90682; // @[Mux.scala 31:69:@36678.4]
  wire [15:0] _T_90683; // @[Mux.scala 31:69:@36679.4]
  wire [15:0] _T_90684; // @[Mux.scala 31:69:@36680.4]
  wire [15:0] _T_90685; // @[Mux.scala 31:69:@36681.4]
  wire [15:0] _T_90686; // @[Mux.scala 31:69:@36682.4]
  wire [15:0] _T_90687; // @[Mux.scala 31:69:@36683.4]
  wire  _T_90688; // @[OneHot.scala 66:30:@36684.4]
  wire  _T_90689; // @[OneHot.scala 66:30:@36685.4]
  wire  _T_90690; // @[OneHot.scala 66:30:@36686.4]
  wire  _T_90691; // @[OneHot.scala 66:30:@36687.4]
  wire  _T_90692; // @[OneHot.scala 66:30:@36688.4]
  wire  _T_90693; // @[OneHot.scala 66:30:@36689.4]
  wire  _T_90694; // @[OneHot.scala 66:30:@36690.4]
  wire  _T_90695; // @[OneHot.scala 66:30:@36691.4]
  wire  _T_90696; // @[OneHot.scala 66:30:@36692.4]
  wire  _T_90697; // @[OneHot.scala 66:30:@36693.4]
  wire  _T_90698; // @[OneHot.scala 66:30:@36694.4]
  wire  _T_90699; // @[OneHot.scala 66:30:@36695.4]
  wire  _T_90700; // @[OneHot.scala 66:30:@36696.4]
  wire  _T_90701; // @[OneHot.scala 66:30:@36697.4]
  wire  _T_90702; // @[OneHot.scala 66:30:@36698.4]
  wire  _T_90703; // @[OneHot.scala 66:30:@36699.4]
  wire [15:0] _T_90744; // @[Mux.scala 31:69:@36717.4]
  wire [15:0] _T_90745; // @[Mux.scala 31:69:@36718.4]
  wire [15:0] _T_90746; // @[Mux.scala 31:69:@36719.4]
  wire [15:0] _T_90747; // @[Mux.scala 31:69:@36720.4]
  wire [15:0] _T_90748; // @[Mux.scala 31:69:@36721.4]
  wire [15:0] _T_90749; // @[Mux.scala 31:69:@36722.4]
  wire [15:0] _T_90750; // @[Mux.scala 31:69:@36723.4]
  wire [15:0] _T_90751; // @[Mux.scala 31:69:@36724.4]
  wire [15:0] _T_90752; // @[Mux.scala 31:69:@36725.4]
  wire [15:0] _T_90753; // @[Mux.scala 31:69:@36726.4]
  wire [15:0] _T_90754; // @[Mux.scala 31:69:@36727.4]
  wire [15:0] _T_90755; // @[Mux.scala 31:69:@36728.4]
  wire [15:0] _T_90756; // @[Mux.scala 31:69:@36729.4]
  wire [15:0] _T_90757; // @[Mux.scala 31:69:@36730.4]
  wire [15:0] _T_90758; // @[Mux.scala 31:69:@36731.4]
  wire [15:0] _T_90759; // @[Mux.scala 31:69:@36732.4]
  wire  _T_90760; // @[OneHot.scala 66:30:@36733.4]
  wire  _T_90761; // @[OneHot.scala 66:30:@36734.4]
  wire  _T_90762; // @[OneHot.scala 66:30:@36735.4]
  wire  _T_90763; // @[OneHot.scala 66:30:@36736.4]
  wire  _T_90764; // @[OneHot.scala 66:30:@36737.4]
  wire  _T_90765; // @[OneHot.scala 66:30:@36738.4]
  wire  _T_90766; // @[OneHot.scala 66:30:@36739.4]
  wire  _T_90767; // @[OneHot.scala 66:30:@36740.4]
  wire  _T_90768; // @[OneHot.scala 66:30:@36741.4]
  wire  _T_90769; // @[OneHot.scala 66:30:@36742.4]
  wire  _T_90770; // @[OneHot.scala 66:30:@36743.4]
  wire  _T_90771; // @[OneHot.scala 66:30:@36744.4]
  wire  _T_90772; // @[OneHot.scala 66:30:@36745.4]
  wire  _T_90773; // @[OneHot.scala 66:30:@36746.4]
  wire  _T_90774; // @[OneHot.scala 66:30:@36747.4]
  wire  _T_90775; // @[OneHot.scala 66:30:@36748.4]
  wire [15:0] _T_90816; // @[Mux.scala 31:69:@36766.4]
  wire [15:0] _T_90817; // @[Mux.scala 31:69:@36767.4]
  wire [15:0] _T_90818; // @[Mux.scala 31:69:@36768.4]
  wire [15:0] _T_90819; // @[Mux.scala 31:69:@36769.4]
  wire [15:0] _T_90820; // @[Mux.scala 31:69:@36770.4]
  wire [15:0] _T_90821; // @[Mux.scala 31:69:@36771.4]
  wire [15:0] _T_90822; // @[Mux.scala 31:69:@36772.4]
  wire [15:0] _T_90823; // @[Mux.scala 31:69:@36773.4]
  wire [15:0] _T_90824; // @[Mux.scala 31:69:@36774.4]
  wire [15:0] _T_90825; // @[Mux.scala 31:69:@36775.4]
  wire [15:0] _T_90826; // @[Mux.scala 31:69:@36776.4]
  wire [15:0] _T_90827; // @[Mux.scala 31:69:@36777.4]
  wire [15:0] _T_90828; // @[Mux.scala 31:69:@36778.4]
  wire [15:0] _T_90829; // @[Mux.scala 31:69:@36779.4]
  wire [15:0] _T_90830; // @[Mux.scala 31:69:@36780.4]
  wire [15:0] _T_90831; // @[Mux.scala 31:69:@36781.4]
  wire  _T_90832; // @[OneHot.scala 66:30:@36782.4]
  wire  _T_90833; // @[OneHot.scala 66:30:@36783.4]
  wire  _T_90834; // @[OneHot.scala 66:30:@36784.4]
  wire  _T_90835; // @[OneHot.scala 66:30:@36785.4]
  wire  _T_90836; // @[OneHot.scala 66:30:@36786.4]
  wire  _T_90837; // @[OneHot.scala 66:30:@36787.4]
  wire  _T_90838; // @[OneHot.scala 66:30:@36788.4]
  wire  _T_90839; // @[OneHot.scala 66:30:@36789.4]
  wire  _T_90840; // @[OneHot.scala 66:30:@36790.4]
  wire  _T_90841; // @[OneHot.scala 66:30:@36791.4]
  wire  _T_90842; // @[OneHot.scala 66:30:@36792.4]
  wire  _T_90843; // @[OneHot.scala 66:30:@36793.4]
  wire  _T_90844; // @[OneHot.scala 66:30:@36794.4]
  wire  _T_90845; // @[OneHot.scala 66:30:@36795.4]
  wire  _T_90846; // @[OneHot.scala 66:30:@36796.4]
  wire  _T_90847; // @[OneHot.scala 66:30:@36797.4]
  wire [15:0] _T_90888; // @[Mux.scala 31:69:@36815.4]
  wire [15:0] _T_90889; // @[Mux.scala 31:69:@36816.4]
  wire [15:0] _T_90890; // @[Mux.scala 31:69:@36817.4]
  wire [15:0] _T_90891; // @[Mux.scala 31:69:@36818.4]
  wire [15:0] _T_90892; // @[Mux.scala 31:69:@36819.4]
  wire [15:0] _T_90893; // @[Mux.scala 31:69:@36820.4]
  wire [15:0] _T_90894; // @[Mux.scala 31:69:@36821.4]
  wire [15:0] _T_90895; // @[Mux.scala 31:69:@36822.4]
  wire [15:0] _T_90896; // @[Mux.scala 31:69:@36823.4]
  wire [15:0] _T_90897; // @[Mux.scala 31:69:@36824.4]
  wire [15:0] _T_90898; // @[Mux.scala 31:69:@36825.4]
  wire [15:0] _T_90899; // @[Mux.scala 31:69:@36826.4]
  wire [15:0] _T_90900; // @[Mux.scala 31:69:@36827.4]
  wire [15:0] _T_90901; // @[Mux.scala 31:69:@36828.4]
  wire [15:0] _T_90902; // @[Mux.scala 31:69:@36829.4]
  wire [15:0] _T_90903; // @[Mux.scala 31:69:@36830.4]
  wire  _T_90904; // @[OneHot.scala 66:30:@36831.4]
  wire  _T_90905; // @[OneHot.scala 66:30:@36832.4]
  wire  _T_90906; // @[OneHot.scala 66:30:@36833.4]
  wire  _T_90907; // @[OneHot.scala 66:30:@36834.4]
  wire  _T_90908; // @[OneHot.scala 66:30:@36835.4]
  wire  _T_90909; // @[OneHot.scala 66:30:@36836.4]
  wire  _T_90910; // @[OneHot.scala 66:30:@36837.4]
  wire  _T_90911; // @[OneHot.scala 66:30:@36838.4]
  wire  _T_90912; // @[OneHot.scala 66:30:@36839.4]
  wire  _T_90913; // @[OneHot.scala 66:30:@36840.4]
  wire  _T_90914; // @[OneHot.scala 66:30:@36841.4]
  wire  _T_90915; // @[OneHot.scala 66:30:@36842.4]
  wire  _T_90916; // @[OneHot.scala 66:30:@36843.4]
  wire  _T_90917; // @[OneHot.scala 66:30:@36844.4]
  wire  _T_90918; // @[OneHot.scala 66:30:@36845.4]
  wire  _T_90919; // @[OneHot.scala 66:30:@36846.4]
  wire [15:0] _T_90960; // @[Mux.scala 31:69:@36864.4]
  wire [15:0] _T_90961; // @[Mux.scala 31:69:@36865.4]
  wire [15:0] _T_90962; // @[Mux.scala 31:69:@36866.4]
  wire [15:0] _T_90963; // @[Mux.scala 31:69:@36867.4]
  wire [15:0] _T_90964; // @[Mux.scala 31:69:@36868.4]
  wire [15:0] _T_90965; // @[Mux.scala 31:69:@36869.4]
  wire [15:0] _T_90966; // @[Mux.scala 31:69:@36870.4]
  wire [15:0] _T_90967; // @[Mux.scala 31:69:@36871.4]
  wire [15:0] _T_90968; // @[Mux.scala 31:69:@36872.4]
  wire [15:0] _T_90969; // @[Mux.scala 31:69:@36873.4]
  wire [15:0] _T_90970; // @[Mux.scala 31:69:@36874.4]
  wire [15:0] _T_90971; // @[Mux.scala 31:69:@36875.4]
  wire [15:0] _T_90972; // @[Mux.scala 31:69:@36876.4]
  wire [15:0] _T_90973; // @[Mux.scala 31:69:@36877.4]
  wire [15:0] _T_90974; // @[Mux.scala 31:69:@36878.4]
  wire [15:0] _T_90975; // @[Mux.scala 31:69:@36879.4]
  wire  _T_90976; // @[OneHot.scala 66:30:@36880.4]
  wire  _T_90977; // @[OneHot.scala 66:30:@36881.4]
  wire  _T_90978; // @[OneHot.scala 66:30:@36882.4]
  wire  _T_90979; // @[OneHot.scala 66:30:@36883.4]
  wire  _T_90980; // @[OneHot.scala 66:30:@36884.4]
  wire  _T_90981; // @[OneHot.scala 66:30:@36885.4]
  wire  _T_90982; // @[OneHot.scala 66:30:@36886.4]
  wire  _T_90983; // @[OneHot.scala 66:30:@36887.4]
  wire  _T_90984; // @[OneHot.scala 66:30:@36888.4]
  wire  _T_90985; // @[OneHot.scala 66:30:@36889.4]
  wire  _T_90986; // @[OneHot.scala 66:30:@36890.4]
  wire  _T_90987; // @[OneHot.scala 66:30:@36891.4]
  wire  _T_90988; // @[OneHot.scala 66:30:@36892.4]
  wire  _T_90989; // @[OneHot.scala 66:30:@36893.4]
  wire  _T_90990; // @[OneHot.scala 66:30:@36894.4]
  wire  _T_90991; // @[OneHot.scala 66:30:@36895.4]
  wire [15:0] _T_91032; // @[Mux.scala 31:69:@36913.4]
  wire [15:0] _T_91033; // @[Mux.scala 31:69:@36914.4]
  wire [15:0] _T_91034; // @[Mux.scala 31:69:@36915.4]
  wire [15:0] _T_91035; // @[Mux.scala 31:69:@36916.4]
  wire [15:0] _T_91036; // @[Mux.scala 31:69:@36917.4]
  wire [15:0] _T_91037; // @[Mux.scala 31:69:@36918.4]
  wire [15:0] _T_91038; // @[Mux.scala 31:69:@36919.4]
  wire [15:0] _T_91039; // @[Mux.scala 31:69:@36920.4]
  wire [15:0] _T_91040; // @[Mux.scala 31:69:@36921.4]
  wire [15:0] _T_91041; // @[Mux.scala 31:69:@36922.4]
  wire [15:0] _T_91042; // @[Mux.scala 31:69:@36923.4]
  wire [15:0] _T_91043; // @[Mux.scala 31:69:@36924.4]
  wire [15:0] _T_91044; // @[Mux.scala 31:69:@36925.4]
  wire [15:0] _T_91045; // @[Mux.scala 31:69:@36926.4]
  wire [15:0] _T_91046; // @[Mux.scala 31:69:@36927.4]
  wire [15:0] _T_91047; // @[Mux.scala 31:69:@36928.4]
  wire  _T_91048; // @[OneHot.scala 66:30:@36929.4]
  wire  _T_91049; // @[OneHot.scala 66:30:@36930.4]
  wire  _T_91050; // @[OneHot.scala 66:30:@36931.4]
  wire  _T_91051; // @[OneHot.scala 66:30:@36932.4]
  wire  _T_91052; // @[OneHot.scala 66:30:@36933.4]
  wire  _T_91053; // @[OneHot.scala 66:30:@36934.4]
  wire  _T_91054; // @[OneHot.scala 66:30:@36935.4]
  wire  _T_91055; // @[OneHot.scala 66:30:@36936.4]
  wire  _T_91056; // @[OneHot.scala 66:30:@36937.4]
  wire  _T_91057; // @[OneHot.scala 66:30:@36938.4]
  wire  _T_91058; // @[OneHot.scala 66:30:@36939.4]
  wire  _T_91059; // @[OneHot.scala 66:30:@36940.4]
  wire  _T_91060; // @[OneHot.scala 66:30:@36941.4]
  wire  _T_91061; // @[OneHot.scala 66:30:@36942.4]
  wire  _T_91062; // @[OneHot.scala 66:30:@36943.4]
  wire  _T_91063; // @[OneHot.scala 66:30:@36944.4]
  wire [15:0] _T_91104; // @[Mux.scala 31:69:@36962.4]
  wire [15:0] _T_91105; // @[Mux.scala 31:69:@36963.4]
  wire [15:0] _T_91106; // @[Mux.scala 31:69:@36964.4]
  wire [15:0] _T_91107; // @[Mux.scala 31:69:@36965.4]
  wire [15:0] _T_91108; // @[Mux.scala 31:69:@36966.4]
  wire [15:0] _T_91109; // @[Mux.scala 31:69:@36967.4]
  wire [15:0] _T_91110; // @[Mux.scala 31:69:@36968.4]
  wire [15:0] _T_91111; // @[Mux.scala 31:69:@36969.4]
  wire [15:0] _T_91112; // @[Mux.scala 31:69:@36970.4]
  wire [15:0] _T_91113; // @[Mux.scala 31:69:@36971.4]
  wire [15:0] _T_91114; // @[Mux.scala 31:69:@36972.4]
  wire [15:0] _T_91115; // @[Mux.scala 31:69:@36973.4]
  wire [15:0] _T_91116; // @[Mux.scala 31:69:@36974.4]
  wire [15:0] _T_91117; // @[Mux.scala 31:69:@36975.4]
  wire [15:0] _T_91118; // @[Mux.scala 31:69:@36976.4]
  wire [15:0] _T_91119; // @[Mux.scala 31:69:@36977.4]
  wire  _T_91120; // @[OneHot.scala 66:30:@36978.4]
  wire  _T_91121; // @[OneHot.scala 66:30:@36979.4]
  wire  _T_91122; // @[OneHot.scala 66:30:@36980.4]
  wire  _T_91123; // @[OneHot.scala 66:30:@36981.4]
  wire  _T_91124; // @[OneHot.scala 66:30:@36982.4]
  wire  _T_91125; // @[OneHot.scala 66:30:@36983.4]
  wire  _T_91126; // @[OneHot.scala 66:30:@36984.4]
  wire  _T_91127; // @[OneHot.scala 66:30:@36985.4]
  wire  _T_91128; // @[OneHot.scala 66:30:@36986.4]
  wire  _T_91129; // @[OneHot.scala 66:30:@36987.4]
  wire  _T_91130; // @[OneHot.scala 66:30:@36988.4]
  wire  _T_91131; // @[OneHot.scala 66:30:@36989.4]
  wire  _T_91132; // @[OneHot.scala 66:30:@36990.4]
  wire  _T_91133; // @[OneHot.scala 66:30:@36991.4]
  wire  _T_91134; // @[OneHot.scala 66:30:@36992.4]
  wire  _T_91135; // @[OneHot.scala 66:30:@36993.4]
  wire [15:0] _T_91176; // @[Mux.scala 31:69:@37011.4]
  wire [15:0] _T_91177; // @[Mux.scala 31:69:@37012.4]
  wire [15:0] _T_91178; // @[Mux.scala 31:69:@37013.4]
  wire [15:0] _T_91179; // @[Mux.scala 31:69:@37014.4]
  wire [15:0] _T_91180; // @[Mux.scala 31:69:@37015.4]
  wire [15:0] _T_91181; // @[Mux.scala 31:69:@37016.4]
  wire [15:0] _T_91182; // @[Mux.scala 31:69:@37017.4]
  wire [15:0] _T_91183; // @[Mux.scala 31:69:@37018.4]
  wire [15:0] _T_91184; // @[Mux.scala 31:69:@37019.4]
  wire [15:0] _T_91185; // @[Mux.scala 31:69:@37020.4]
  wire [15:0] _T_91186; // @[Mux.scala 31:69:@37021.4]
  wire [15:0] _T_91187; // @[Mux.scala 31:69:@37022.4]
  wire [15:0] _T_91188; // @[Mux.scala 31:69:@37023.4]
  wire [15:0] _T_91189; // @[Mux.scala 31:69:@37024.4]
  wire [15:0] _T_91190; // @[Mux.scala 31:69:@37025.4]
  wire [15:0] _T_91191; // @[Mux.scala 31:69:@37026.4]
  wire  _T_91192; // @[OneHot.scala 66:30:@37027.4]
  wire  _T_91193; // @[OneHot.scala 66:30:@37028.4]
  wire  _T_91194; // @[OneHot.scala 66:30:@37029.4]
  wire  _T_91195; // @[OneHot.scala 66:30:@37030.4]
  wire  _T_91196; // @[OneHot.scala 66:30:@37031.4]
  wire  _T_91197; // @[OneHot.scala 66:30:@37032.4]
  wire  _T_91198; // @[OneHot.scala 66:30:@37033.4]
  wire  _T_91199; // @[OneHot.scala 66:30:@37034.4]
  wire  _T_91200; // @[OneHot.scala 66:30:@37035.4]
  wire  _T_91201; // @[OneHot.scala 66:30:@37036.4]
  wire  _T_91202; // @[OneHot.scala 66:30:@37037.4]
  wire  _T_91203; // @[OneHot.scala 66:30:@37038.4]
  wire  _T_91204; // @[OneHot.scala 66:30:@37039.4]
  wire  _T_91205; // @[OneHot.scala 66:30:@37040.4]
  wire  _T_91206; // @[OneHot.scala 66:30:@37041.4]
  wire  _T_91207; // @[OneHot.scala 66:30:@37042.4]
  wire [15:0] _T_91248; // @[Mux.scala 31:69:@37060.4]
  wire [15:0] _T_91249; // @[Mux.scala 31:69:@37061.4]
  wire [15:0] _T_91250; // @[Mux.scala 31:69:@37062.4]
  wire [15:0] _T_91251; // @[Mux.scala 31:69:@37063.4]
  wire [15:0] _T_91252; // @[Mux.scala 31:69:@37064.4]
  wire [15:0] _T_91253; // @[Mux.scala 31:69:@37065.4]
  wire [15:0] _T_91254; // @[Mux.scala 31:69:@37066.4]
  wire [15:0] _T_91255; // @[Mux.scala 31:69:@37067.4]
  wire [15:0] _T_91256; // @[Mux.scala 31:69:@37068.4]
  wire [15:0] _T_91257; // @[Mux.scala 31:69:@37069.4]
  wire [15:0] _T_91258; // @[Mux.scala 31:69:@37070.4]
  wire [15:0] _T_91259; // @[Mux.scala 31:69:@37071.4]
  wire [15:0] _T_91260; // @[Mux.scala 31:69:@37072.4]
  wire [15:0] _T_91261; // @[Mux.scala 31:69:@37073.4]
  wire [15:0] _T_91262; // @[Mux.scala 31:69:@37074.4]
  wire [15:0] _T_91263; // @[Mux.scala 31:69:@37075.4]
  wire  _T_91264; // @[OneHot.scala 66:30:@37076.4]
  wire  _T_91265; // @[OneHot.scala 66:30:@37077.4]
  wire  _T_91266; // @[OneHot.scala 66:30:@37078.4]
  wire  _T_91267; // @[OneHot.scala 66:30:@37079.4]
  wire  _T_91268; // @[OneHot.scala 66:30:@37080.4]
  wire  _T_91269; // @[OneHot.scala 66:30:@37081.4]
  wire  _T_91270; // @[OneHot.scala 66:30:@37082.4]
  wire  _T_91271; // @[OneHot.scala 66:30:@37083.4]
  wire  _T_91272; // @[OneHot.scala 66:30:@37084.4]
  wire  _T_91273; // @[OneHot.scala 66:30:@37085.4]
  wire  _T_91274; // @[OneHot.scala 66:30:@37086.4]
  wire  _T_91275; // @[OneHot.scala 66:30:@37087.4]
  wire  _T_91276; // @[OneHot.scala 66:30:@37088.4]
  wire  _T_91277; // @[OneHot.scala 66:30:@37089.4]
  wire  _T_91278; // @[OneHot.scala 66:30:@37090.4]
  wire  _T_91279; // @[OneHot.scala 66:30:@37091.4]
  wire [15:0] _T_91320; // @[Mux.scala 31:69:@37109.4]
  wire [15:0] _T_91321; // @[Mux.scala 31:69:@37110.4]
  wire [15:0] _T_91322; // @[Mux.scala 31:69:@37111.4]
  wire [15:0] _T_91323; // @[Mux.scala 31:69:@37112.4]
  wire [15:0] _T_91324; // @[Mux.scala 31:69:@37113.4]
  wire [15:0] _T_91325; // @[Mux.scala 31:69:@37114.4]
  wire [15:0] _T_91326; // @[Mux.scala 31:69:@37115.4]
  wire [15:0] _T_91327; // @[Mux.scala 31:69:@37116.4]
  wire [15:0] _T_91328; // @[Mux.scala 31:69:@37117.4]
  wire [15:0] _T_91329; // @[Mux.scala 31:69:@37118.4]
  wire [15:0] _T_91330; // @[Mux.scala 31:69:@37119.4]
  wire [15:0] _T_91331; // @[Mux.scala 31:69:@37120.4]
  wire [15:0] _T_91332; // @[Mux.scala 31:69:@37121.4]
  wire [15:0] _T_91333; // @[Mux.scala 31:69:@37122.4]
  wire [15:0] _T_91334; // @[Mux.scala 31:69:@37123.4]
  wire [15:0] _T_91335; // @[Mux.scala 31:69:@37124.4]
  wire  _T_91336; // @[OneHot.scala 66:30:@37125.4]
  wire  _T_91337; // @[OneHot.scala 66:30:@37126.4]
  wire  _T_91338; // @[OneHot.scala 66:30:@37127.4]
  wire  _T_91339; // @[OneHot.scala 66:30:@37128.4]
  wire  _T_91340; // @[OneHot.scala 66:30:@37129.4]
  wire  _T_91341; // @[OneHot.scala 66:30:@37130.4]
  wire  _T_91342; // @[OneHot.scala 66:30:@37131.4]
  wire  _T_91343; // @[OneHot.scala 66:30:@37132.4]
  wire  _T_91344; // @[OneHot.scala 66:30:@37133.4]
  wire  _T_91345; // @[OneHot.scala 66:30:@37134.4]
  wire  _T_91346; // @[OneHot.scala 66:30:@37135.4]
  wire  _T_91347; // @[OneHot.scala 66:30:@37136.4]
  wire  _T_91348; // @[OneHot.scala 66:30:@37137.4]
  wire  _T_91349; // @[OneHot.scala 66:30:@37138.4]
  wire  _T_91350; // @[OneHot.scala 66:30:@37139.4]
  wire  _T_91351; // @[OneHot.scala 66:30:@37140.4]
  wire [15:0] _T_91392; // @[Mux.scala 31:69:@37158.4]
  wire [15:0] _T_91393; // @[Mux.scala 31:69:@37159.4]
  wire [15:0] _T_91394; // @[Mux.scala 31:69:@37160.4]
  wire [15:0] _T_91395; // @[Mux.scala 31:69:@37161.4]
  wire [15:0] _T_91396; // @[Mux.scala 31:69:@37162.4]
  wire [15:0] _T_91397; // @[Mux.scala 31:69:@37163.4]
  wire [15:0] _T_91398; // @[Mux.scala 31:69:@37164.4]
  wire [15:0] _T_91399; // @[Mux.scala 31:69:@37165.4]
  wire [15:0] _T_91400; // @[Mux.scala 31:69:@37166.4]
  wire [15:0] _T_91401; // @[Mux.scala 31:69:@37167.4]
  wire [15:0] _T_91402; // @[Mux.scala 31:69:@37168.4]
  wire [15:0] _T_91403; // @[Mux.scala 31:69:@37169.4]
  wire [15:0] _T_91404; // @[Mux.scala 31:69:@37170.4]
  wire [15:0] _T_91405; // @[Mux.scala 31:69:@37171.4]
  wire [15:0] _T_91406; // @[Mux.scala 31:69:@37172.4]
  wire [15:0] _T_91407; // @[Mux.scala 31:69:@37173.4]
  wire  _T_91408; // @[OneHot.scala 66:30:@37174.4]
  wire  _T_91409; // @[OneHot.scala 66:30:@37175.4]
  wire  _T_91410; // @[OneHot.scala 66:30:@37176.4]
  wire  _T_91411; // @[OneHot.scala 66:30:@37177.4]
  wire  _T_91412; // @[OneHot.scala 66:30:@37178.4]
  wire  _T_91413; // @[OneHot.scala 66:30:@37179.4]
  wire  _T_91414; // @[OneHot.scala 66:30:@37180.4]
  wire  _T_91415; // @[OneHot.scala 66:30:@37181.4]
  wire  _T_91416; // @[OneHot.scala 66:30:@37182.4]
  wire  _T_91417; // @[OneHot.scala 66:30:@37183.4]
  wire  _T_91418; // @[OneHot.scala 66:30:@37184.4]
  wire  _T_91419; // @[OneHot.scala 66:30:@37185.4]
  wire  _T_91420; // @[OneHot.scala 66:30:@37186.4]
  wire  _T_91421; // @[OneHot.scala 66:30:@37187.4]
  wire  _T_91422; // @[OneHot.scala 66:30:@37188.4]
  wire  _T_91423; // @[OneHot.scala 66:30:@37189.4]
  wire [15:0] _T_91464; // @[Mux.scala 31:69:@37207.4]
  wire [15:0] _T_91465; // @[Mux.scala 31:69:@37208.4]
  wire [15:0] _T_91466; // @[Mux.scala 31:69:@37209.4]
  wire [15:0] _T_91467; // @[Mux.scala 31:69:@37210.4]
  wire [15:0] _T_91468; // @[Mux.scala 31:69:@37211.4]
  wire [15:0] _T_91469; // @[Mux.scala 31:69:@37212.4]
  wire [15:0] _T_91470; // @[Mux.scala 31:69:@37213.4]
  wire [15:0] _T_91471; // @[Mux.scala 31:69:@37214.4]
  wire [15:0] _T_91472; // @[Mux.scala 31:69:@37215.4]
  wire [15:0] _T_91473; // @[Mux.scala 31:69:@37216.4]
  wire [15:0] _T_91474; // @[Mux.scala 31:69:@37217.4]
  wire [15:0] _T_91475; // @[Mux.scala 31:69:@37218.4]
  wire [15:0] _T_91476; // @[Mux.scala 31:69:@37219.4]
  wire [15:0] _T_91477; // @[Mux.scala 31:69:@37220.4]
  wire [15:0] _T_91478; // @[Mux.scala 31:69:@37221.4]
  wire [15:0] _T_91479; // @[Mux.scala 31:69:@37222.4]
  wire  _T_91480; // @[OneHot.scala 66:30:@37223.4]
  wire  _T_91481; // @[OneHot.scala 66:30:@37224.4]
  wire  _T_91482; // @[OneHot.scala 66:30:@37225.4]
  wire  _T_91483; // @[OneHot.scala 66:30:@37226.4]
  wire  _T_91484; // @[OneHot.scala 66:30:@37227.4]
  wire  _T_91485; // @[OneHot.scala 66:30:@37228.4]
  wire  _T_91486; // @[OneHot.scala 66:30:@37229.4]
  wire  _T_91487; // @[OneHot.scala 66:30:@37230.4]
  wire  _T_91488; // @[OneHot.scala 66:30:@37231.4]
  wire  _T_91489; // @[OneHot.scala 66:30:@37232.4]
  wire  _T_91490; // @[OneHot.scala 66:30:@37233.4]
  wire  _T_91491; // @[OneHot.scala 66:30:@37234.4]
  wire  _T_91492; // @[OneHot.scala 66:30:@37235.4]
  wire  _T_91493; // @[OneHot.scala 66:30:@37236.4]
  wire  _T_91494; // @[OneHot.scala 66:30:@37237.4]
  wire  _T_91495; // @[OneHot.scala 66:30:@37238.4]
  wire [15:0] _T_91536; // @[Mux.scala 31:69:@37256.4]
  wire [15:0] _T_91537; // @[Mux.scala 31:69:@37257.4]
  wire [15:0] _T_91538; // @[Mux.scala 31:69:@37258.4]
  wire [15:0] _T_91539; // @[Mux.scala 31:69:@37259.4]
  wire [15:0] _T_91540; // @[Mux.scala 31:69:@37260.4]
  wire [15:0] _T_91541; // @[Mux.scala 31:69:@37261.4]
  wire [15:0] _T_91542; // @[Mux.scala 31:69:@37262.4]
  wire [15:0] _T_91543; // @[Mux.scala 31:69:@37263.4]
  wire [15:0] _T_91544; // @[Mux.scala 31:69:@37264.4]
  wire [15:0] _T_91545; // @[Mux.scala 31:69:@37265.4]
  wire [15:0] _T_91546; // @[Mux.scala 31:69:@37266.4]
  wire [15:0] _T_91547; // @[Mux.scala 31:69:@37267.4]
  wire [15:0] _T_91548; // @[Mux.scala 31:69:@37268.4]
  wire [15:0] _T_91549; // @[Mux.scala 31:69:@37269.4]
  wire [15:0] _T_91550; // @[Mux.scala 31:69:@37270.4]
  wire [15:0] _T_91551; // @[Mux.scala 31:69:@37271.4]
  wire  _T_91552; // @[OneHot.scala 66:30:@37272.4]
  wire  _T_91553; // @[OneHot.scala 66:30:@37273.4]
  wire  _T_91554; // @[OneHot.scala 66:30:@37274.4]
  wire  _T_91555; // @[OneHot.scala 66:30:@37275.4]
  wire  _T_91556; // @[OneHot.scala 66:30:@37276.4]
  wire  _T_91557; // @[OneHot.scala 66:30:@37277.4]
  wire  _T_91558; // @[OneHot.scala 66:30:@37278.4]
  wire  _T_91559; // @[OneHot.scala 66:30:@37279.4]
  wire  _T_91560; // @[OneHot.scala 66:30:@37280.4]
  wire  _T_91561; // @[OneHot.scala 66:30:@37281.4]
  wire  _T_91562; // @[OneHot.scala 66:30:@37282.4]
  wire  _T_91563; // @[OneHot.scala 66:30:@37283.4]
  wire  _T_91564; // @[OneHot.scala 66:30:@37284.4]
  wire  _T_91565; // @[OneHot.scala 66:30:@37285.4]
  wire  _T_91566; // @[OneHot.scala 66:30:@37286.4]
  wire  _T_91567; // @[OneHot.scala 66:30:@37287.4]
  wire [7:0] _T_91632; // @[Mux.scala 19:72:@37311.4]
  wire [15:0] _T_91640; // @[Mux.scala 19:72:@37319.4]
  wire [15:0] _T_91642; // @[Mux.scala 19:72:@37320.4]
  wire [7:0] _T_91649; // @[Mux.scala 19:72:@37327.4]
  wire [15:0] _T_91657; // @[Mux.scala 19:72:@37335.4]
  wire [15:0] _T_91659; // @[Mux.scala 19:72:@37336.4]
  wire [7:0] _T_91666; // @[Mux.scala 19:72:@37343.4]
  wire [15:0] _T_91674; // @[Mux.scala 19:72:@37351.4]
  wire [15:0] _T_91676; // @[Mux.scala 19:72:@37352.4]
  wire [7:0] _T_91683; // @[Mux.scala 19:72:@37359.4]
  wire [15:0] _T_91691; // @[Mux.scala 19:72:@37367.4]
  wire [15:0] _T_91693; // @[Mux.scala 19:72:@37368.4]
  wire [7:0] _T_91700; // @[Mux.scala 19:72:@37375.4]
  wire [15:0] _T_91708; // @[Mux.scala 19:72:@37383.4]
  wire [15:0] _T_91710; // @[Mux.scala 19:72:@37384.4]
  wire [7:0] _T_91717; // @[Mux.scala 19:72:@37391.4]
  wire [15:0] _T_91725; // @[Mux.scala 19:72:@37399.4]
  wire [15:0] _T_91727; // @[Mux.scala 19:72:@37400.4]
  wire [7:0] _T_91734; // @[Mux.scala 19:72:@37407.4]
  wire [15:0] _T_91742; // @[Mux.scala 19:72:@37415.4]
  wire [15:0] _T_91744; // @[Mux.scala 19:72:@37416.4]
  wire [7:0] _T_91751; // @[Mux.scala 19:72:@37423.4]
  wire [15:0] _T_91759; // @[Mux.scala 19:72:@37431.4]
  wire [15:0] _T_91761; // @[Mux.scala 19:72:@37432.4]
  wire [7:0] _T_91768; // @[Mux.scala 19:72:@37439.4]
  wire [15:0] _T_91776; // @[Mux.scala 19:72:@37447.4]
  wire [15:0] _T_91778; // @[Mux.scala 19:72:@37448.4]
  wire [7:0] _T_91785; // @[Mux.scala 19:72:@37455.4]
  wire [15:0] _T_91793; // @[Mux.scala 19:72:@37463.4]
  wire [15:0] _T_91795; // @[Mux.scala 19:72:@37464.4]
  wire [7:0] _T_91802; // @[Mux.scala 19:72:@37471.4]
  wire [15:0] _T_91810; // @[Mux.scala 19:72:@37479.4]
  wire [15:0] _T_91812; // @[Mux.scala 19:72:@37480.4]
  wire [7:0] _T_91819; // @[Mux.scala 19:72:@37487.4]
  wire [15:0] _T_91827; // @[Mux.scala 19:72:@37495.4]
  wire [15:0] _T_91829; // @[Mux.scala 19:72:@37496.4]
  wire [7:0] _T_91836; // @[Mux.scala 19:72:@37503.4]
  wire [15:0] _T_91844; // @[Mux.scala 19:72:@37511.4]
  wire [15:0] _T_91846; // @[Mux.scala 19:72:@37512.4]
  wire [7:0] _T_91853; // @[Mux.scala 19:72:@37519.4]
  wire [15:0] _T_91861; // @[Mux.scala 19:72:@37527.4]
  wire [15:0] _T_91863; // @[Mux.scala 19:72:@37528.4]
  wire [7:0] _T_91870; // @[Mux.scala 19:72:@37535.4]
  wire [15:0] _T_91878; // @[Mux.scala 19:72:@37543.4]
  wire [15:0] _T_91880; // @[Mux.scala 19:72:@37544.4]
  wire [7:0] _T_91887; // @[Mux.scala 19:72:@37551.4]
  wire [15:0] _T_91895; // @[Mux.scala 19:72:@37559.4]
  wire [15:0] _T_91897; // @[Mux.scala 19:72:@37560.4]
  wire [15:0] _T_91898; // @[Mux.scala 19:72:@37561.4]
  wire [15:0] _T_91899; // @[Mux.scala 19:72:@37562.4]
  wire [15:0] _T_91900; // @[Mux.scala 19:72:@37563.4]
  wire [15:0] _T_91901; // @[Mux.scala 19:72:@37564.4]
  wire [15:0] _T_91902; // @[Mux.scala 19:72:@37565.4]
  wire [15:0] _T_91903; // @[Mux.scala 19:72:@37566.4]
  wire [15:0] _T_91904; // @[Mux.scala 19:72:@37567.4]
  wire [15:0] _T_91905; // @[Mux.scala 19:72:@37568.4]
  wire [15:0] _T_91906; // @[Mux.scala 19:72:@37569.4]
  wire [15:0] _T_91907; // @[Mux.scala 19:72:@37570.4]
  wire [15:0] _T_91908; // @[Mux.scala 19:72:@37571.4]
  wire [15:0] _T_91909; // @[Mux.scala 19:72:@37572.4]
  wire [15:0] _T_91910; // @[Mux.scala 19:72:@37573.4]
  wire [15:0] _T_91911; // @[Mux.scala 19:72:@37574.4]
  wire [15:0] _T_91912; // @[Mux.scala 19:72:@37575.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@37579.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@37581.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@37583.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@37585.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@37587.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@37589.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@37591.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@37593.4]
  wire  priorityLoadRequest_8; // @[Mux.scala 19:72:@37595.4]
  wire  priorityLoadRequest_9; // @[Mux.scala 19:72:@37597.4]
  wire  priorityLoadRequest_10; // @[Mux.scala 19:72:@37599.4]
  wire  priorityLoadRequest_11; // @[Mux.scala 19:72:@37601.4]
  wire  priorityLoadRequest_12; // @[Mux.scala 19:72:@37603.4]
  wire  priorityLoadRequest_13; // @[Mux.scala 19:72:@37605.4]
  wire  priorityLoadRequest_14; // @[Mux.scala 19:72:@37607.4]
  wire  priorityLoadRequest_15; // @[Mux.scala 19:72:@37609.4]
  wire  _GEN_1920; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1921; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1922; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1923; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1924; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1925; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1926; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1927; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1928; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1929; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1930; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1931; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1932; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1933; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1934; // @[LoadQueue.scala 208:31:@37629.4]
  wire  _GEN_1935; // @[LoadQueue.scala 208:31:@37629.4]
  wire [7:0] _T_92307; // @[LoadQueue.scala 238:58:@37847.8]
  wire [15:0] _T_92315; // @[LoadQueue.scala 238:58:@37855.8]
  wire [7:0] _T_92322; // @[LoadQueue.scala 238:96:@37862.8]
  wire [15:0] _T_92330; // @[LoadQueue.scala 238:96:@37870.8]
  wire  _T_92331; // @[LoadQueue.scala 238:61:@37871.8]
  wire  _T_92332; // @[LoadQueue.scala 237:64:@37872.8]
  wire  _GEN_1969; // @[LoadQueue.scala 230:110:@37804.6]
  wire  bypassRequest_0; // @[LoadQueue.scala 229:71:@37798.4]
  wire  _GEN_1936; // @[LoadQueue.scala 217:34:@37686.6]
  wire  _GEN_1937; // @[LoadQueue.scala 215:23:@37682.4]
  wire [7:0] _T_92391; // @[LoadQueue.scala 238:58:@37929.8]
  wire [15:0] _T_92399; // @[LoadQueue.scala 238:58:@37937.8]
  wire [7:0] _T_92406; // @[LoadQueue.scala 238:96:@37944.8]
  wire [15:0] _T_92414; // @[LoadQueue.scala 238:96:@37952.8]
  wire  _T_92415; // @[LoadQueue.scala 238:61:@37953.8]
  wire  _T_92416; // @[LoadQueue.scala 237:64:@37954.8]
  wire  _GEN_1973; // @[LoadQueue.scala 230:110:@37886.6]
  wire  bypassRequest_1; // @[LoadQueue.scala 229:71:@37880.4]
  wire  _GEN_1938; // @[LoadQueue.scala 217:34:@37693.6]
  wire  _GEN_1939; // @[LoadQueue.scala 215:23:@37689.4]
  wire [7:0] _T_92475; // @[LoadQueue.scala 238:58:@38011.8]
  wire [15:0] _T_92483; // @[LoadQueue.scala 238:58:@38019.8]
  wire [7:0] _T_92490; // @[LoadQueue.scala 238:96:@38026.8]
  wire [15:0] _T_92498; // @[LoadQueue.scala 238:96:@38034.8]
  wire  _T_92499; // @[LoadQueue.scala 238:61:@38035.8]
  wire  _T_92500; // @[LoadQueue.scala 237:64:@38036.8]
  wire  _GEN_1977; // @[LoadQueue.scala 230:110:@37968.6]
  wire  bypassRequest_2; // @[LoadQueue.scala 229:71:@37962.4]
  wire  _GEN_1940; // @[LoadQueue.scala 217:34:@37700.6]
  wire  _GEN_1941; // @[LoadQueue.scala 215:23:@37696.4]
  wire [7:0] _T_92559; // @[LoadQueue.scala 238:58:@38093.8]
  wire [15:0] _T_92567; // @[LoadQueue.scala 238:58:@38101.8]
  wire [7:0] _T_92574; // @[LoadQueue.scala 238:96:@38108.8]
  wire [15:0] _T_92582; // @[LoadQueue.scala 238:96:@38116.8]
  wire  _T_92583; // @[LoadQueue.scala 238:61:@38117.8]
  wire  _T_92584; // @[LoadQueue.scala 237:64:@38118.8]
  wire  _GEN_1981; // @[LoadQueue.scala 230:110:@38050.6]
  wire  bypassRequest_3; // @[LoadQueue.scala 229:71:@38044.4]
  wire  _GEN_1942; // @[LoadQueue.scala 217:34:@37707.6]
  wire  _GEN_1943; // @[LoadQueue.scala 215:23:@37703.4]
  wire [7:0] _T_92643; // @[LoadQueue.scala 238:58:@38175.8]
  wire [15:0] _T_92651; // @[LoadQueue.scala 238:58:@38183.8]
  wire [7:0] _T_92658; // @[LoadQueue.scala 238:96:@38190.8]
  wire [15:0] _T_92666; // @[LoadQueue.scala 238:96:@38198.8]
  wire  _T_92667; // @[LoadQueue.scala 238:61:@38199.8]
  wire  _T_92668; // @[LoadQueue.scala 237:64:@38200.8]
  wire  _GEN_1985; // @[LoadQueue.scala 230:110:@38132.6]
  wire  bypassRequest_4; // @[LoadQueue.scala 229:71:@38126.4]
  wire  _GEN_1944; // @[LoadQueue.scala 217:34:@37714.6]
  wire  _GEN_1945; // @[LoadQueue.scala 215:23:@37710.4]
  wire [7:0] _T_92727; // @[LoadQueue.scala 238:58:@38257.8]
  wire [15:0] _T_92735; // @[LoadQueue.scala 238:58:@38265.8]
  wire [7:0] _T_92742; // @[LoadQueue.scala 238:96:@38272.8]
  wire [15:0] _T_92750; // @[LoadQueue.scala 238:96:@38280.8]
  wire  _T_92751; // @[LoadQueue.scala 238:61:@38281.8]
  wire  _T_92752; // @[LoadQueue.scala 237:64:@38282.8]
  wire  _GEN_1989; // @[LoadQueue.scala 230:110:@38214.6]
  wire  bypassRequest_5; // @[LoadQueue.scala 229:71:@38208.4]
  wire  _GEN_1946; // @[LoadQueue.scala 217:34:@37721.6]
  wire  _GEN_1947; // @[LoadQueue.scala 215:23:@37717.4]
  wire [7:0] _T_92811; // @[LoadQueue.scala 238:58:@38339.8]
  wire [15:0] _T_92819; // @[LoadQueue.scala 238:58:@38347.8]
  wire [7:0] _T_92826; // @[LoadQueue.scala 238:96:@38354.8]
  wire [15:0] _T_92834; // @[LoadQueue.scala 238:96:@38362.8]
  wire  _T_92835; // @[LoadQueue.scala 238:61:@38363.8]
  wire  _T_92836; // @[LoadQueue.scala 237:64:@38364.8]
  wire  _GEN_1993; // @[LoadQueue.scala 230:110:@38296.6]
  wire  bypassRequest_6; // @[LoadQueue.scala 229:71:@38290.4]
  wire  _GEN_1948; // @[LoadQueue.scala 217:34:@37728.6]
  wire  _GEN_1949; // @[LoadQueue.scala 215:23:@37724.4]
  wire [7:0] _T_92895; // @[LoadQueue.scala 238:58:@38421.8]
  wire [15:0] _T_92903; // @[LoadQueue.scala 238:58:@38429.8]
  wire [7:0] _T_92910; // @[LoadQueue.scala 238:96:@38436.8]
  wire [15:0] _T_92918; // @[LoadQueue.scala 238:96:@38444.8]
  wire  _T_92919; // @[LoadQueue.scala 238:61:@38445.8]
  wire  _T_92920; // @[LoadQueue.scala 237:64:@38446.8]
  wire  _GEN_1997; // @[LoadQueue.scala 230:110:@38378.6]
  wire  bypassRequest_7; // @[LoadQueue.scala 229:71:@38372.4]
  wire  _GEN_1950; // @[LoadQueue.scala 217:34:@37735.6]
  wire  _GEN_1951; // @[LoadQueue.scala 215:23:@37731.4]
  wire [7:0] _T_92979; // @[LoadQueue.scala 238:58:@38503.8]
  wire [15:0] _T_92987; // @[LoadQueue.scala 238:58:@38511.8]
  wire [7:0] _T_92994; // @[LoadQueue.scala 238:96:@38518.8]
  wire [15:0] _T_93002; // @[LoadQueue.scala 238:96:@38526.8]
  wire  _T_93003; // @[LoadQueue.scala 238:61:@38527.8]
  wire  _T_93004; // @[LoadQueue.scala 237:64:@38528.8]
  wire  _GEN_2001; // @[LoadQueue.scala 230:110:@38460.6]
  wire  bypassRequest_8; // @[LoadQueue.scala 229:71:@38454.4]
  wire  _GEN_1952; // @[LoadQueue.scala 217:34:@37742.6]
  wire  _GEN_1953; // @[LoadQueue.scala 215:23:@37738.4]
  wire [7:0] _T_93063; // @[LoadQueue.scala 238:58:@38585.8]
  wire [15:0] _T_93071; // @[LoadQueue.scala 238:58:@38593.8]
  wire [7:0] _T_93078; // @[LoadQueue.scala 238:96:@38600.8]
  wire [15:0] _T_93086; // @[LoadQueue.scala 238:96:@38608.8]
  wire  _T_93087; // @[LoadQueue.scala 238:61:@38609.8]
  wire  _T_93088; // @[LoadQueue.scala 237:64:@38610.8]
  wire  _GEN_2005; // @[LoadQueue.scala 230:110:@38542.6]
  wire  bypassRequest_9; // @[LoadQueue.scala 229:71:@38536.4]
  wire  _GEN_1954; // @[LoadQueue.scala 217:34:@37749.6]
  wire  _GEN_1955; // @[LoadQueue.scala 215:23:@37745.4]
  wire [7:0] _T_93147; // @[LoadQueue.scala 238:58:@38667.8]
  wire [15:0] _T_93155; // @[LoadQueue.scala 238:58:@38675.8]
  wire [7:0] _T_93162; // @[LoadQueue.scala 238:96:@38682.8]
  wire [15:0] _T_93170; // @[LoadQueue.scala 238:96:@38690.8]
  wire  _T_93171; // @[LoadQueue.scala 238:61:@38691.8]
  wire  _T_93172; // @[LoadQueue.scala 237:64:@38692.8]
  wire  _GEN_2009; // @[LoadQueue.scala 230:110:@38624.6]
  wire  bypassRequest_10; // @[LoadQueue.scala 229:71:@38618.4]
  wire  _GEN_1956; // @[LoadQueue.scala 217:34:@37756.6]
  wire  _GEN_1957; // @[LoadQueue.scala 215:23:@37752.4]
  wire [7:0] _T_93231; // @[LoadQueue.scala 238:58:@38749.8]
  wire [15:0] _T_93239; // @[LoadQueue.scala 238:58:@38757.8]
  wire [7:0] _T_93246; // @[LoadQueue.scala 238:96:@38764.8]
  wire [15:0] _T_93254; // @[LoadQueue.scala 238:96:@38772.8]
  wire  _T_93255; // @[LoadQueue.scala 238:61:@38773.8]
  wire  _T_93256; // @[LoadQueue.scala 237:64:@38774.8]
  wire  _GEN_2013; // @[LoadQueue.scala 230:110:@38706.6]
  wire  bypassRequest_11; // @[LoadQueue.scala 229:71:@38700.4]
  wire  _GEN_1958; // @[LoadQueue.scala 217:34:@37763.6]
  wire  _GEN_1959; // @[LoadQueue.scala 215:23:@37759.4]
  wire [7:0] _T_93315; // @[LoadQueue.scala 238:58:@38831.8]
  wire [15:0] _T_93323; // @[LoadQueue.scala 238:58:@38839.8]
  wire [7:0] _T_93330; // @[LoadQueue.scala 238:96:@38846.8]
  wire [15:0] _T_93338; // @[LoadQueue.scala 238:96:@38854.8]
  wire  _T_93339; // @[LoadQueue.scala 238:61:@38855.8]
  wire  _T_93340; // @[LoadQueue.scala 237:64:@38856.8]
  wire  _GEN_2017; // @[LoadQueue.scala 230:110:@38788.6]
  wire  bypassRequest_12; // @[LoadQueue.scala 229:71:@38782.4]
  wire  _GEN_1960; // @[LoadQueue.scala 217:34:@37770.6]
  wire  _GEN_1961; // @[LoadQueue.scala 215:23:@37766.4]
  wire [7:0] _T_93399; // @[LoadQueue.scala 238:58:@38913.8]
  wire [15:0] _T_93407; // @[LoadQueue.scala 238:58:@38921.8]
  wire [7:0] _T_93414; // @[LoadQueue.scala 238:96:@38928.8]
  wire [15:0] _T_93422; // @[LoadQueue.scala 238:96:@38936.8]
  wire  _T_93423; // @[LoadQueue.scala 238:61:@38937.8]
  wire  _T_93424; // @[LoadQueue.scala 237:64:@38938.8]
  wire  _GEN_2021; // @[LoadQueue.scala 230:110:@38870.6]
  wire  bypassRequest_13; // @[LoadQueue.scala 229:71:@38864.4]
  wire  _GEN_1962; // @[LoadQueue.scala 217:34:@37777.6]
  wire  _GEN_1963; // @[LoadQueue.scala 215:23:@37773.4]
  wire [7:0] _T_93483; // @[LoadQueue.scala 238:58:@38995.8]
  wire [15:0] _T_93491; // @[LoadQueue.scala 238:58:@39003.8]
  wire [7:0] _T_93498; // @[LoadQueue.scala 238:96:@39010.8]
  wire [15:0] _T_93506; // @[LoadQueue.scala 238:96:@39018.8]
  wire  _T_93507; // @[LoadQueue.scala 238:61:@39019.8]
  wire  _T_93508; // @[LoadQueue.scala 237:64:@39020.8]
  wire  _GEN_2025; // @[LoadQueue.scala 230:110:@38952.6]
  wire  bypassRequest_14; // @[LoadQueue.scala 229:71:@38946.4]
  wire  _GEN_1964; // @[LoadQueue.scala 217:34:@37784.6]
  wire  _GEN_1965; // @[LoadQueue.scala 215:23:@37780.4]
  wire [7:0] _T_93567; // @[LoadQueue.scala 238:58:@39077.8]
  wire [15:0] _T_93575; // @[LoadQueue.scala 238:58:@39085.8]
  wire [7:0] _T_93582; // @[LoadQueue.scala 238:96:@39092.8]
  wire [15:0] _T_93590; // @[LoadQueue.scala 238:96:@39100.8]
  wire  _T_93591; // @[LoadQueue.scala 238:61:@39101.8]
  wire  _T_93592; // @[LoadQueue.scala 237:64:@39102.8]
  wire  _GEN_2029; // @[LoadQueue.scala 230:110:@39034.6]
  wire  bypassRequest_15; // @[LoadQueue.scala 229:71:@39028.4]
  wire  _GEN_1966; // @[LoadQueue.scala 217:34:@37791.6]
  wire  _GEN_1967; // @[LoadQueue.scala 215:23:@37787.4]
  wire  _T_93596; // @[LoadQueue.scala 247:28:@39108.4]
  wire  _T_93597; // @[LoadQueue.scala 247:28:@39109.4]
  wire  _T_93598; // @[LoadQueue.scala 247:28:@39110.4]
  wire  _T_93599; // @[LoadQueue.scala 247:28:@39111.4]
  wire  _T_93600; // @[LoadQueue.scala 247:28:@39112.4]
  wire  _T_93601; // @[LoadQueue.scala 247:28:@39113.4]
  wire  _T_93602; // @[LoadQueue.scala 247:28:@39114.4]
  wire  _T_93603; // @[LoadQueue.scala 247:28:@39115.4]
  wire  _T_93604; // @[LoadQueue.scala 247:28:@39116.4]
  wire  _T_93605; // @[LoadQueue.scala 247:28:@39117.4]
  wire  _T_93606; // @[LoadQueue.scala 247:28:@39118.4]
  wire  _T_93607; // @[LoadQueue.scala 247:28:@39119.4]
  wire  _T_93608; // @[LoadQueue.scala 247:28:@39120.4]
  wire  _T_93609; // @[LoadQueue.scala 247:28:@39121.4]
  wire  _T_93610; // @[LoadQueue.scala 247:28:@39122.4]
  wire [3:0] _T_93627; // @[Mux.scala 31:69:@39124.6]
  wire [3:0] _T_93628; // @[Mux.scala 31:69:@39125.6]
  wire [3:0] _T_93629; // @[Mux.scala 31:69:@39126.6]
  wire [3:0] _T_93630; // @[Mux.scala 31:69:@39127.6]
  wire [3:0] _T_93631; // @[Mux.scala 31:69:@39128.6]
  wire [3:0] _T_93632; // @[Mux.scala 31:69:@39129.6]
  wire [3:0] _T_93633; // @[Mux.scala 31:69:@39130.6]
  wire [3:0] _T_93634; // @[Mux.scala 31:69:@39131.6]
  wire [3:0] _T_93635; // @[Mux.scala 31:69:@39132.6]
  wire [3:0] _T_93636; // @[Mux.scala 31:69:@39133.6]
  wire [3:0] _T_93637; // @[Mux.scala 31:69:@39134.6]
  wire [3:0] _T_93638; // @[Mux.scala 31:69:@39135.6]
  wire [3:0] _T_93639; // @[Mux.scala 31:69:@39136.6]
  wire [3:0] _T_93640; // @[Mux.scala 31:69:@39137.6]
  wire [3:0] _T_93641; // @[Mux.scala 31:69:@39138.6]
  wire [31:0] _GEN_2033; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2034; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2035; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2036; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2037; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2038; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2039; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2040; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2041; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2042; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2043; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2044; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2045; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2046; // @[LoadQueue.scala 248:24:@39139.6]
  wire [31:0] _GEN_2047; // @[LoadQueue.scala 248:24:@39139.6]
  wire  _T_93649; // @[LoadQueue.scala 261:41:@39150.6]
  wire  _GEN_2050; // @[LoadQueue.scala 261:62:@39151.6]
  wire  _GEN_2051; // @[LoadQueue.scala 259:25:@39146.4]
  wire  _T_93652; // @[LoadQueue.scala 261:41:@39158.6]
  wire  _GEN_2052; // @[LoadQueue.scala 261:62:@39159.6]
  wire  _GEN_2053; // @[LoadQueue.scala 259:25:@39154.4]
  wire  _T_93655; // @[LoadQueue.scala 261:41:@39166.6]
  wire  _GEN_2054; // @[LoadQueue.scala 261:62:@39167.6]
  wire  _GEN_2055; // @[LoadQueue.scala 259:25:@39162.4]
  wire  _T_93658; // @[LoadQueue.scala 261:41:@39174.6]
  wire  _GEN_2056; // @[LoadQueue.scala 261:62:@39175.6]
  wire  _GEN_2057; // @[LoadQueue.scala 259:25:@39170.4]
  wire  _T_93661; // @[LoadQueue.scala 261:41:@39182.6]
  wire  _GEN_2058; // @[LoadQueue.scala 261:62:@39183.6]
  wire  _GEN_2059; // @[LoadQueue.scala 259:25:@39178.4]
  wire  _T_93664; // @[LoadQueue.scala 261:41:@39190.6]
  wire  _GEN_2060; // @[LoadQueue.scala 261:62:@39191.6]
  wire  _GEN_2061; // @[LoadQueue.scala 259:25:@39186.4]
  wire  _T_93667; // @[LoadQueue.scala 261:41:@39198.6]
  wire  _GEN_2062; // @[LoadQueue.scala 261:62:@39199.6]
  wire  _GEN_2063; // @[LoadQueue.scala 259:25:@39194.4]
  wire  _T_93670; // @[LoadQueue.scala 261:41:@39206.6]
  wire  _GEN_2064; // @[LoadQueue.scala 261:62:@39207.6]
  wire  _GEN_2065; // @[LoadQueue.scala 259:25:@39202.4]
  wire  _T_93673; // @[LoadQueue.scala 261:41:@39214.6]
  wire  _GEN_2066; // @[LoadQueue.scala 261:62:@39215.6]
  wire  _GEN_2067; // @[LoadQueue.scala 259:25:@39210.4]
  wire  _T_93676; // @[LoadQueue.scala 261:41:@39222.6]
  wire  _GEN_2068; // @[LoadQueue.scala 261:62:@39223.6]
  wire  _GEN_2069; // @[LoadQueue.scala 259:25:@39218.4]
  wire  _T_93679; // @[LoadQueue.scala 261:41:@39230.6]
  wire  _GEN_2070; // @[LoadQueue.scala 261:62:@39231.6]
  wire  _GEN_2071; // @[LoadQueue.scala 259:25:@39226.4]
  wire  _T_93682; // @[LoadQueue.scala 261:41:@39238.6]
  wire  _GEN_2072; // @[LoadQueue.scala 261:62:@39239.6]
  wire  _GEN_2073; // @[LoadQueue.scala 259:25:@39234.4]
  wire  _T_93685; // @[LoadQueue.scala 261:41:@39246.6]
  wire  _GEN_2074; // @[LoadQueue.scala 261:62:@39247.6]
  wire  _GEN_2075; // @[LoadQueue.scala 259:25:@39242.4]
  wire  _T_93688; // @[LoadQueue.scala 261:41:@39254.6]
  wire  _GEN_2076; // @[LoadQueue.scala 261:62:@39255.6]
  wire  _GEN_2077; // @[LoadQueue.scala 259:25:@39250.4]
  wire  _T_93691; // @[LoadQueue.scala 261:41:@39262.6]
  wire  _GEN_2078; // @[LoadQueue.scala 261:62:@39263.6]
  wire  _GEN_2079; // @[LoadQueue.scala 259:25:@39258.4]
  wire  _T_93694; // @[LoadQueue.scala 261:41:@39270.6]
  wire  _GEN_2080; // @[LoadQueue.scala 261:62:@39271.6]
  wire  _GEN_2081; // @[LoadQueue.scala 259:25:@39266.4]
  wire [31:0] _GEN_2082; // @[LoadQueue.scala 269:44:@39278.6]
  wire [31:0] _GEN_2083; // @[LoadQueue.scala 267:32:@39274.4]
  wire [31:0] _GEN_2084; // @[LoadQueue.scala 269:44:@39285.6]
  wire [31:0] _GEN_2085; // @[LoadQueue.scala 267:32:@39281.4]
  wire [31:0] _GEN_2086; // @[LoadQueue.scala 269:44:@39292.6]
  wire [31:0] _GEN_2087; // @[LoadQueue.scala 267:32:@39288.4]
  wire [31:0] _GEN_2088; // @[LoadQueue.scala 269:44:@39299.6]
  wire [31:0] _GEN_2089; // @[LoadQueue.scala 267:32:@39295.4]
  wire [31:0] _GEN_2090; // @[LoadQueue.scala 269:44:@39306.6]
  wire [31:0] _GEN_2091; // @[LoadQueue.scala 267:32:@39302.4]
  wire [31:0] _GEN_2092; // @[LoadQueue.scala 269:44:@39313.6]
  wire [31:0] _GEN_2093; // @[LoadQueue.scala 267:32:@39309.4]
  wire [31:0] _GEN_2094; // @[LoadQueue.scala 269:44:@39320.6]
  wire [31:0] _GEN_2095; // @[LoadQueue.scala 267:32:@39316.4]
  wire [31:0] _GEN_2096; // @[LoadQueue.scala 269:44:@39327.6]
  wire [31:0] _GEN_2097; // @[LoadQueue.scala 267:32:@39323.4]
  wire [31:0] _GEN_2098; // @[LoadQueue.scala 269:44:@39334.6]
  wire [31:0] _GEN_2099; // @[LoadQueue.scala 267:32:@39330.4]
  wire [31:0] _GEN_2100; // @[LoadQueue.scala 269:44:@39341.6]
  wire [31:0] _GEN_2101; // @[LoadQueue.scala 267:32:@39337.4]
  wire [31:0] _GEN_2102; // @[LoadQueue.scala 269:44:@39348.6]
  wire [31:0] _GEN_2103; // @[LoadQueue.scala 267:32:@39344.4]
  wire [31:0] _GEN_2104; // @[LoadQueue.scala 269:44:@39355.6]
  wire [31:0] _GEN_2105; // @[LoadQueue.scala 267:32:@39351.4]
  wire [31:0] _GEN_2106; // @[LoadQueue.scala 269:44:@39362.6]
  wire [31:0] _GEN_2107; // @[LoadQueue.scala 267:32:@39358.4]
  wire [31:0] _GEN_2108; // @[LoadQueue.scala 269:44:@39369.6]
  wire [31:0] _GEN_2109; // @[LoadQueue.scala 267:32:@39365.4]
  wire [31:0] _GEN_2110; // @[LoadQueue.scala 269:44:@39376.6]
  wire [31:0] _GEN_2111; // @[LoadQueue.scala 267:32:@39372.4]
  wire [31:0] _GEN_2112; // @[LoadQueue.scala 269:44:@39383.6]
  wire [31:0] _GEN_2113; // @[LoadQueue.scala 267:32:@39379.4]
  wire  entriesPorts_0_0; // @[LoadQueue.scala 286:69:@39387.4]
  wire  entriesPorts_0_1; // @[LoadQueue.scala 286:69:@39389.4]
  wire  entriesPorts_0_2; // @[LoadQueue.scala 286:69:@39391.4]
  wire  entriesPorts_0_3; // @[LoadQueue.scala 286:69:@39393.4]
  wire  entriesPorts_0_4; // @[LoadQueue.scala 286:69:@39395.4]
  wire  entriesPorts_0_5; // @[LoadQueue.scala 286:69:@39397.4]
  wire  entriesPorts_0_6; // @[LoadQueue.scala 286:69:@39399.4]
  wire  entriesPorts_0_7; // @[LoadQueue.scala 286:69:@39401.4]
  wire  entriesPorts_0_8; // @[LoadQueue.scala 286:69:@39403.4]
  wire  entriesPorts_0_9; // @[LoadQueue.scala 286:69:@39405.4]
  wire  entriesPorts_0_10; // @[LoadQueue.scala 286:69:@39407.4]
  wire  entriesPorts_0_11; // @[LoadQueue.scala 286:69:@39409.4]
  wire  entriesPorts_0_12; // @[LoadQueue.scala 286:69:@39411.4]
  wire  entriesPorts_0_13; // @[LoadQueue.scala 286:69:@39413.4]
  wire  entriesPorts_0_14; // @[LoadQueue.scala 286:69:@39415.4]
  wire  entriesPorts_0_15; // @[LoadQueue.scala 286:69:@39417.4]
  wire  _T_94179; // @[LoadQueue.scala 298:86:@39421.4]
  wire  _T_94180; // @[LoadQueue.scala 298:83:@39422.4]
  wire  _T_94182; // @[LoadQueue.scala 298:86:@39423.4]
  wire  _T_94183; // @[LoadQueue.scala 298:83:@39424.4]
  wire  _T_94185; // @[LoadQueue.scala 298:86:@39425.4]
  wire  _T_94186; // @[LoadQueue.scala 298:83:@39426.4]
  wire  _T_94188; // @[LoadQueue.scala 298:86:@39427.4]
  wire  _T_94189; // @[LoadQueue.scala 298:83:@39428.4]
  wire  _T_94191; // @[LoadQueue.scala 298:86:@39429.4]
  wire  _T_94192; // @[LoadQueue.scala 298:83:@39430.4]
  wire  _T_94194; // @[LoadQueue.scala 298:86:@39431.4]
  wire  _T_94195; // @[LoadQueue.scala 298:83:@39432.4]
  wire  _T_94197; // @[LoadQueue.scala 298:86:@39433.4]
  wire  _T_94198; // @[LoadQueue.scala 298:83:@39434.4]
  wire  _T_94200; // @[LoadQueue.scala 298:86:@39435.4]
  wire  _T_94201; // @[LoadQueue.scala 298:83:@39436.4]
  wire  _T_94203; // @[LoadQueue.scala 298:86:@39437.4]
  wire  _T_94204; // @[LoadQueue.scala 298:83:@39438.4]
  wire  _T_94206; // @[LoadQueue.scala 298:86:@39439.4]
  wire  _T_94207; // @[LoadQueue.scala 298:83:@39440.4]
  wire  _T_94209; // @[LoadQueue.scala 298:86:@39441.4]
  wire  _T_94210; // @[LoadQueue.scala 298:83:@39442.4]
  wire  _T_94212; // @[LoadQueue.scala 298:86:@39443.4]
  wire  _T_94213; // @[LoadQueue.scala 298:83:@39444.4]
  wire  _T_94215; // @[LoadQueue.scala 298:86:@39445.4]
  wire  _T_94216; // @[LoadQueue.scala 298:83:@39446.4]
  wire  _T_94218; // @[LoadQueue.scala 298:86:@39447.4]
  wire  _T_94219; // @[LoadQueue.scala 298:83:@39448.4]
  wire  _T_94221; // @[LoadQueue.scala 298:86:@39449.4]
  wire  _T_94222; // @[LoadQueue.scala 298:83:@39450.4]
  wire  _T_94224; // @[LoadQueue.scala 298:86:@39451.4]
  wire  _T_94225; // @[LoadQueue.scala 298:83:@39452.4]
  wire [15:0] _T_94308; // @[Mux.scala 31:69:@39506.4]
  wire [15:0] _T_94309; // @[Mux.scala 31:69:@39507.4]
  wire [15:0] _T_94310; // @[Mux.scala 31:69:@39508.4]
  wire [15:0] _T_94311; // @[Mux.scala 31:69:@39509.4]
  wire [15:0] _T_94312; // @[Mux.scala 31:69:@39510.4]
  wire [15:0] _T_94313; // @[Mux.scala 31:69:@39511.4]
  wire [15:0] _T_94314; // @[Mux.scala 31:69:@39512.4]
  wire [15:0] _T_94315; // @[Mux.scala 31:69:@39513.4]
  wire [15:0] _T_94316; // @[Mux.scala 31:69:@39514.4]
  wire [15:0] _T_94317; // @[Mux.scala 31:69:@39515.4]
  wire [15:0] _T_94318; // @[Mux.scala 31:69:@39516.4]
  wire [15:0] _T_94319; // @[Mux.scala 31:69:@39517.4]
  wire [15:0] _T_94320; // @[Mux.scala 31:69:@39518.4]
  wire [15:0] _T_94321; // @[Mux.scala 31:69:@39519.4]
  wire [15:0] _T_94322; // @[Mux.scala 31:69:@39520.4]
  wire [15:0] _T_94323; // @[Mux.scala 31:69:@39521.4]
  wire  _T_94324; // @[OneHot.scala 66:30:@39522.4]
  wire  _T_94325; // @[OneHot.scala 66:30:@39523.4]
  wire  _T_94326; // @[OneHot.scala 66:30:@39524.4]
  wire  _T_94327; // @[OneHot.scala 66:30:@39525.4]
  wire  _T_94328; // @[OneHot.scala 66:30:@39526.4]
  wire  _T_94329; // @[OneHot.scala 66:30:@39527.4]
  wire  _T_94330; // @[OneHot.scala 66:30:@39528.4]
  wire  _T_94331; // @[OneHot.scala 66:30:@39529.4]
  wire  _T_94332; // @[OneHot.scala 66:30:@39530.4]
  wire  _T_94333; // @[OneHot.scala 66:30:@39531.4]
  wire  _T_94334; // @[OneHot.scala 66:30:@39532.4]
  wire  _T_94335; // @[OneHot.scala 66:30:@39533.4]
  wire  _T_94336; // @[OneHot.scala 66:30:@39534.4]
  wire  _T_94337; // @[OneHot.scala 66:30:@39535.4]
  wire  _T_94338; // @[OneHot.scala 66:30:@39536.4]
  wire  _T_94339; // @[OneHot.scala 66:30:@39537.4]
  wire [15:0] _T_94380; // @[Mux.scala 31:69:@39555.4]
  wire [15:0] _T_94381; // @[Mux.scala 31:69:@39556.4]
  wire [15:0] _T_94382; // @[Mux.scala 31:69:@39557.4]
  wire [15:0] _T_94383; // @[Mux.scala 31:69:@39558.4]
  wire [15:0] _T_94384; // @[Mux.scala 31:69:@39559.4]
  wire [15:0] _T_94385; // @[Mux.scala 31:69:@39560.4]
  wire [15:0] _T_94386; // @[Mux.scala 31:69:@39561.4]
  wire [15:0] _T_94387; // @[Mux.scala 31:69:@39562.4]
  wire [15:0] _T_94388; // @[Mux.scala 31:69:@39563.4]
  wire [15:0] _T_94389; // @[Mux.scala 31:69:@39564.4]
  wire [15:0] _T_94390; // @[Mux.scala 31:69:@39565.4]
  wire [15:0] _T_94391; // @[Mux.scala 31:69:@39566.4]
  wire [15:0] _T_94392; // @[Mux.scala 31:69:@39567.4]
  wire [15:0] _T_94393; // @[Mux.scala 31:69:@39568.4]
  wire [15:0] _T_94394; // @[Mux.scala 31:69:@39569.4]
  wire [15:0] _T_94395; // @[Mux.scala 31:69:@39570.4]
  wire  _T_94396; // @[OneHot.scala 66:30:@39571.4]
  wire  _T_94397; // @[OneHot.scala 66:30:@39572.4]
  wire  _T_94398; // @[OneHot.scala 66:30:@39573.4]
  wire  _T_94399; // @[OneHot.scala 66:30:@39574.4]
  wire  _T_94400; // @[OneHot.scala 66:30:@39575.4]
  wire  _T_94401; // @[OneHot.scala 66:30:@39576.4]
  wire  _T_94402; // @[OneHot.scala 66:30:@39577.4]
  wire  _T_94403; // @[OneHot.scala 66:30:@39578.4]
  wire  _T_94404; // @[OneHot.scala 66:30:@39579.4]
  wire  _T_94405; // @[OneHot.scala 66:30:@39580.4]
  wire  _T_94406; // @[OneHot.scala 66:30:@39581.4]
  wire  _T_94407; // @[OneHot.scala 66:30:@39582.4]
  wire  _T_94408; // @[OneHot.scala 66:30:@39583.4]
  wire  _T_94409; // @[OneHot.scala 66:30:@39584.4]
  wire  _T_94410; // @[OneHot.scala 66:30:@39585.4]
  wire  _T_94411; // @[OneHot.scala 66:30:@39586.4]
  wire [15:0] _T_94452; // @[Mux.scala 31:69:@39604.4]
  wire [15:0] _T_94453; // @[Mux.scala 31:69:@39605.4]
  wire [15:0] _T_94454; // @[Mux.scala 31:69:@39606.4]
  wire [15:0] _T_94455; // @[Mux.scala 31:69:@39607.4]
  wire [15:0] _T_94456; // @[Mux.scala 31:69:@39608.4]
  wire [15:0] _T_94457; // @[Mux.scala 31:69:@39609.4]
  wire [15:0] _T_94458; // @[Mux.scala 31:69:@39610.4]
  wire [15:0] _T_94459; // @[Mux.scala 31:69:@39611.4]
  wire [15:0] _T_94460; // @[Mux.scala 31:69:@39612.4]
  wire [15:0] _T_94461; // @[Mux.scala 31:69:@39613.4]
  wire [15:0] _T_94462; // @[Mux.scala 31:69:@39614.4]
  wire [15:0] _T_94463; // @[Mux.scala 31:69:@39615.4]
  wire [15:0] _T_94464; // @[Mux.scala 31:69:@39616.4]
  wire [15:0] _T_94465; // @[Mux.scala 31:69:@39617.4]
  wire [15:0] _T_94466; // @[Mux.scala 31:69:@39618.4]
  wire [15:0] _T_94467; // @[Mux.scala 31:69:@39619.4]
  wire  _T_94468; // @[OneHot.scala 66:30:@39620.4]
  wire  _T_94469; // @[OneHot.scala 66:30:@39621.4]
  wire  _T_94470; // @[OneHot.scala 66:30:@39622.4]
  wire  _T_94471; // @[OneHot.scala 66:30:@39623.4]
  wire  _T_94472; // @[OneHot.scala 66:30:@39624.4]
  wire  _T_94473; // @[OneHot.scala 66:30:@39625.4]
  wire  _T_94474; // @[OneHot.scala 66:30:@39626.4]
  wire  _T_94475; // @[OneHot.scala 66:30:@39627.4]
  wire  _T_94476; // @[OneHot.scala 66:30:@39628.4]
  wire  _T_94477; // @[OneHot.scala 66:30:@39629.4]
  wire  _T_94478; // @[OneHot.scala 66:30:@39630.4]
  wire  _T_94479; // @[OneHot.scala 66:30:@39631.4]
  wire  _T_94480; // @[OneHot.scala 66:30:@39632.4]
  wire  _T_94481; // @[OneHot.scala 66:30:@39633.4]
  wire  _T_94482; // @[OneHot.scala 66:30:@39634.4]
  wire  _T_94483; // @[OneHot.scala 66:30:@39635.4]
  wire [15:0] _T_94524; // @[Mux.scala 31:69:@39653.4]
  wire [15:0] _T_94525; // @[Mux.scala 31:69:@39654.4]
  wire [15:0] _T_94526; // @[Mux.scala 31:69:@39655.4]
  wire [15:0] _T_94527; // @[Mux.scala 31:69:@39656.4]
  wire [15:0] _T_94528; // @[Mux.scala 31:69:@39657.4]
  wire [15:0] _T_94529; // @[Mux.scala 31:69:@39658.4]
  wire [15:0] _T_94530; // @[Mux.scala 31:69:@39659.4]
  wire [15:0] _T_94531; // @[Mux.scala 31:69:@39660.4]
  wire [15:0] _T_94532; // @[Mux.scala 31:69:@39661.4]
  wire [15:0] _T_94533; // @[Mux.scala 31:69:@39662.4]
  wire [15:0] _T_94534; // @[Mux.scala 31:69:@39663.4]
  wire [15:0] _T_94535; // @[Mux.scala 31:69:@39664.4]
  wire [15:0] _T_94536; // @[Mux.scala 31:69:@39665.4]
  wire [15:0] _T_94537; // @[Mux.scala 31:69:@39666.4]
  wire [15:0] _T_94538; // @[Mux.scala 31:69:@39667.4]
  wire [15:0] _T_94539; // @[Mux.scala 31:69:@39668.4]
  wire  _T_94540; // @[OneHot.scala 66:30:@39669.4]
  wire  _T_94541; // @[OneHot.scala 66:30:@39670.4]
  wire  _T_94542; // @[OneHot.scala 66:30:@39671.4]
  wire  _T_94543; // @[OneHot.scala 66:30:@39672.4]
  wire  _T_94544; // @[OneHot.scala 66:30:@39673.4]
  wire  _T_94545; // @[OneHot.scala 66:30:@39674.4]
  wire  _T_94546; // @[OneHot.scala 66:30:@39675.4]
  wire  _T_94547; // @[OneHot.scala 66:30:@39676.4]
  wire  _T_94548; // @[OneHot.scala 66:30:@39677.4]
  wire  _T_94549; // @[OneHot.scala 66:30:@39678.4]
  wire  _T_94550; // @[OneHot.scala 66:30:@39679.4]
  wire  _T_94551; // @[OneHot.scala 66:30:@39680.4]
  wire  _T_94552; // @[OneHot.scala 66:30:@39681.4]
  wire  _T_94553; // @[OneHot.scala 66:30:@39682.4]
  wire  _T_94554; // @[OneHot.scala 66:30:@39683.4]
  wire  _T_94555; // @[OneHot.scala 66:30:@39684.4]
  wire [15:0] _T_94596; // @[Mux.scala 31:69:@39702.4]
  wire [15:0] _T_94597; // @[Mux.scala 31:69:@39703.4]
  wire [15:0] _T_94598; // @[Mux.scala 31:69:@39704.4]
  wire [15:0] _T_94599; // @[Mux.scala 31:69:@39705.4]
  wire [15:0] _T_94600; // @[Mux.scala 31:69:@39706.4]
  wire [15:0] _T_94601; // @[Mux.scala 31:69:@39707.4]
  wire [15:0] _T_94602; // @[Mux.scala 31:69:@39708.4]
  wire [15:0] _T_94603; // @[Mux.scala 31:69:@39709.4]
  wire [15:0] _T_94604; // @[Mux.scala 31:69:@39710.4]
  wire [15:0] _T_94605; // @[Mux.scala 31:69:@39711.4]
  wire [15:0] _T_94606; // @[Mux.scala 31:69:@39712.4]
  wire [15:0] _T_94607; // @[Mux.scala 31:69:@39713.4]
  wire [15:0] _T_94608; // @[Mux.scala 31:69:@39714.4]
  wire [15:0] _T_94609; // @[Mux.scala 31:69:@39715.4]
  wire [15:0] _T_94610; // @[Mux.scala 31:69:@39716.4]
  wire [15:0] _T_94611; // @[Mux.scala 31:69:@39717.4]
  wire  _T_94612; // @[OneHot.scala 66:30:@39718.4]
  wire  _T_94613; // @[OneHot.scala 66:30:@39719.4]
  wire  _T_94614; // @[OneHot.scala 66:30:@39720.4]
  wire  _T_94615; // @[OneHot.scala 66:30:@39721.4]
  wire  _T_94616; // @[OneHot.scala 66:30:@39722.4]
  wire  _T_94617; // @[OneHot.scala 66:30:@39723.4]
  wire  _T_94618; // @[OneHot.scala 66:30:@39724.4]
  wire  _T_94619; // @[OneHot.scala 66:30:@39725.4]
  wire  _T_94620; // @[OneHot.scala 66:30:@39726.4]
  wire  _T_94621; // @[OneHot.scala 66:30:@39727.4]
  wire  _T_94622; // @[OneHot.scala 66:30:@39728.4]
  wire  _T_94623; // @[OneHot.scala 66:30:@39729.4]
  wire  _T_94624; // @[OneHot.scala 66:30:@39730.4]
  wire  _T_94625; // @[OneHot.scala 66:30:@39731.4]
  wire  _T_94626; // @[OneHot.scala 66:30:@39732.4]
  wire  _T_94627; // @[OneHot.scala 66:30:@39733.4]
  wire [15:0] _T_94668; // @[Mux.scala 31:69:@39751.4]
  wire [15:0] _T_94669; // @[Mux.scala 31:69:@39752.4]
  wire [15:0] _T_94670; // @[Mux.scala 31:69:@39753.4]
  wire [15:0] _T_94671; // @[Mux.scala 31:69:@39754.4]
  wire [15:0] _T_94672; // @[Mux.scala 31:69:@39755.4]
  wire [15:0] _T_94673; // @[Mux.scala 31:69:@39756.4]
  wire [15:0] _T_94674; // @[Mux.scala 31:69:@39757.4]
  wire [15:0] _T_94675; // @[Mux.scala 31:69:@39758.4]
  wire [15:0] _T_94676; // @[Mux.scala 31:69:@39759.4]
  wire [15:0] _T_94677; // @[Mux.scala 31:69:@39760.4]
  wire [15:0] _T_94678; // @[Mux.scala 31:69:@39761.4]
  wire [15:0] _T_94679; // @[Mux.scala 31:69:@39762.4]
  wire [15:0] _T_94680; // @[Mux.scala 31:69:@39763.4]
  wire [15:0] _T_94681; // @[Mux.scala 31:69:@39764.4]
  wire [15:0] _T_94682; // @[Mux.scala 31:69:@39765.4]
  wire [15:0] _T_94683; // @[Mux.scala 31:69:@39766.4]
  wire  _T_94684; // @[OneHot.scala 66:30:@39767.4]
  wire  _T_94685; // @[OneHot.scala 66:30:@39768.4]
  wire  _T_94686; // @[OneHot.scala 66:30:@39769.4]
  wire  _T_94687; // @[OneHot.scala 66:30:@39770.4]
  wire  _T_94688; // @[OneHot.scala 66:30:@39771.4]
  wire  _T_94689; // @[OneHot.scala 66:30:@39772.4]
  wire  _T_94690; // @[OneHot.scala 66:30:@39773.4]
  wire  _T_94691; // @[OneHot.scala 66:30:@39774.4]
  wire  _T_94692; // @[OneHot.scala 66:30:@39775.4]
  wire  _T_94693; // @[OneHot.scala 66:30:@39776.4]
  wire  _T_94694; // @[OneHot.scala 66:30:@39777.4]
  wire  _T_94695; // @[OneHot.scala 66:30:@39778.4]
  wire  _T_94696; // @[OneHot.scala 66:30:@39779.4]
  wire  _T_94697; // @[OneHot.scala 66:30:@39780.4]
  wire  _T_94698; // @[OneHot.scala 66:30:@39781.4]
  wire  _T_94699; // @[OneHot.scala 66:30:@39782.4]
  wire [15:0] _T_94740; // @[Mux.scala 31:69:@39800.4]
  wire [15:0] _T_94741; // @[Mux.scala 31:69:@39801.4]
  wire [15:0] _T_94742; // @[Mux.scala 31:69:@39802.4]
  wire [15:0] _T_94743; // @[Mux.scala 31:69:@39803.4]
  wire [15:0] _T_94744; // @[Mux.scala 31:69:@39804.4]
  wire [15:0] _T_94745; // @[Mux.scala 31:69:@39805.4]
  wire [15:0] _T_94746; // @[Mux.scala 31:69:@39806.4]
  wire [15:0] _T_94747; // @[Mux.scala 31:69:@39807.4]
  wire [15:0] _T_94748; // @[Mux.scala 31:69:@39808.4]
  wire [15:0] _T_94749; // @[Mux.scala 31:69:@39809.4]
  wire [15:0] _T_94750; // @[Mux.scala 31:69:@39810.4]
  wire [15:0] _T_94751; // @[Mux.scala 31:69:@39811.4]
  wire [15:0] _T_94752; // @[Mux.scala 31:69:@39812.4]
  wire [15:0] _T_94753; // @[Mux.scala 31:69:@39813.4]
  wire [15:0] _T_94754; // @[Mux.scala 31:69:@39814.4]
  wire [15:0] _T_94755; // @[Mux.scala 31:69:@39815.4]
  wire  _T_94756; // @[OneHot.scala 66:30:@39816.4]
  wire  _T_94757; // @[OneHot.scala 66:30:@39817.4]
  wire  _T_94758; // @[OneHot.scala 66:30:@39818.4]
  wire  _T_94759; // @[OneHot.scala 66:30:@39819.4]
  wire  _T_94760; // @[OneHot.scala 66:30:@39820.4]
  wire  _T_94761; // @[OneHot.scala 66:30:@39821.4]
  wire  _T_94762; // @[OneHot.scala 66:30:@39822.4]
  wire  _T_94763; // @[OneHot.scala 66:30:@39823.4]
  wire  _T_94764; // @[OneHot.scala 66:30:@39824.4]
  wire  _T_94765; // @[OneHot.scala 66:30:@39825.4]
  wire  _T_94766; // @[OneHot.scala 66:30:@39826.4]
  wire  _T_94767; // @[OneHot.scala 66:30:@39827.4]
  wire  _T_94768; // @[OneHot.scala 66:30:@39828.4]
  wire  _T_94769; // @[OneHot.scala 66:30:@39829.4]
  wire  _T_94770; // @[OneHot.scala 66:30:@39830.4]
  wire  _T_94771; // @[OneHot.scala 66:30:@39831.4]
  wire [15:0] _T_94812; // @[Mux.scala 31:69:@39849.4]
  wire [15:0] _T_94813; // @[Mux.scala 31:69:@39850.4]
  wire [15:0] _T_94814; // @[Mux.scala 31:69:@39851.4]
  wire [15:0] _T_94815; // @[Mux.scala 31:69:@39852.4]
  wire [15:0] _T_94816; // @[Mux.scala 31:69:@39853.4]
  wire [15:0] _T_94817; // @[Mux.scala 31:69:@39854.4]
  wire [15:0] _T_94818; // @[Mux.scala 31:69:@39855.4]
  wire [15:0] _T_94819; // @[Mux.scala 31:69:@39856.4]
  wire [15:0] _T_94820; // @[Mux.scala 31:69:@39857.4]
  wire [15:0] _T_94821; // @[Mux.scala 31:69:@39858.4]
  wire [15:0] _T_94822; // @[Mux.scala 31:69:@39859.4]
  wire [15:0] _T_94823; // @[Mux.scala 31:69:@39860.4]
  wire [15:0] _T_94824; // @[Mux.scala 31:69:@39861.4]
  wire [15:0] _T_94825; // @[Mux.scala 31:69:@39862.4]
  wire [15:0] _T_94826; // @[Mux.scala 31:69:@39863.4]
  wire [15:0] _T_94827; // @[Mux.scala 31:69:@39864.4]
  wire  _T_94828; // @[OneHot.scala 66:30:@39865.4]
  wire  _T_94829; // @[OneHot.scala 66:30:@39866.4]
  wire  _T_94830; // @[OneHot.scala 66:30:@39867.4]
  wire  _T_94831; // @[OneHot.scala 66:30:@39868.4]
  wire  _T_94832; // @[OneHot.scala 66:30:@39869.4]
  wire  _T_94833; // @[OneHot.scala 66:30:@39870.4]
  wire  _T_94834; // @[OneHot.scala 66:30:@39871.4]
  wire  _T_94835; // @[OneHot.scala 66:30:@39872.4]
  wire  _T_94836; // @[OneHot.scala 66:30:@39873.4]
  wire  _T_94837; // @[OneHot.scala 66:30:@39874.4]
  wire  _T_94838; // @[OneHot.scala 66:30:@39875.4]
  wire  _T_94839; // @[OneHot.scala 66:30:@39876.4]
  wire  _T_94840; // @[OneHot.scala 66:30:@39877.4]
  wire  _T_94841; // @[OneHot.scala 66:30:@39878.4]
  wire  _T_94842; // @[OneHot.scala 66:30:@39879.4]
  wire  _T_94843; // @[OneHot.scala 66:30:@39880.4]
  wire [15:0] _T_94884; // @[Mux.scala 31:69:@39898.4]
  wire [15:0] _T_94885; // @[Mux.scala 31:69:@39899.4]
  wire [15:0] _T_94886; // @[Mux.scala 31:69:@39900.4]
  wire [15:0] _T_94887; // @[Mux.scala 31:69:@39901.4]
  wire [15:0] _T_94888; // @[Mux.scala 31:69:@39902.4]
  wire [15:0] _T_94889; // @[Mux.scala 31:69:@39903.4]
  wire [15:0] _T_94890; // @[Mux.scala 31:69:@39904.4]
  wire [15:0] _T_94891; // @[Mux.scala 31:69:@39905.4]
  wire [15:0] _T_94892; // @[Mux.scala 31:69:@39906.4]
  wire [15:0] _T_94893; // @[Mux.scala 31:69:@39907.4]
  wire [15:0] _T_94894; // @[Mux.scala 31:69:@39908.4]
  wire [15:0] _T_94895; // @[Mux.scala 31:69:@39909.4]
  wire [15:0] _T_94896; // @[Mux.scala 31:69:@39910.4]
  wire [15:0] _T_94897; // @[Mux.scala 31:69:@39911.4]
  wire [15:0] _T_94898; // @[Mux.scala 31:69:@39912.4]
  wire [15:0] _T_94899; // @[Mux.scala 31:69:@39913.4]
  wire  _T_94900; // @[OneHot.scala 66:30:@39914.4]
  wire  _T_94901; // @[OneHot.scala 66:30:@39915.4]
  wire  _T_94902; // @[OneHot.scala 66:30:@39916.4]
  wire  _T_94903; // @[OneHot.scala 66:30:@39917.4]
  wire  _T_94904; // @[OneHot.scala 66:30:@39918.4]
  wire  _T_94905; // @[OneHot.scala 66:30:@39919.4]
  wire  _T_94906; // @[OneHot.scala 66:30:@39920.4]
  wire  _T_94907; // @[OneHot.scala 66:30:@39921.4]
  wire  _T_94908; // @[OneHot.scala 66:30:@39922.4]
  wire  _T_94909; // @[OneHot.scala 66:30:@39923.4]
  wire  _T_94910; // @[OneHot.scala 66:30:@39924.4]
  wire  _T_94911; // @[OneHot.scala 66:30:@39925.4]
  wire  _T_94912; // @[OneHot.scala 66:30:@39926.4]
  wire  _T_94913; // @[OneHot.scala 66:30:@39927.4]
  wire  _T_94914; // @[OneHot.scala 66:30:@39928.4]
  wire  _T_94915; // @[OneHot.scala 66:30:@39929.4]
  wire [15:0] _T_94956; // @[Mux.scala 31:69:@39947.4]
  wire [15:0] _T_94957; // @[Mux.scala 31:69:@39948.4]
  wire [15:0] _T_94958; // @[Mux.scala 31:69:@39949.4]
  wire [15:0] _T_94959; // @[Mux.scala 31:69:@39950.4]
  wire [15:0] _T_94960; // @[Mux.scala 31:69:@39951.4]
  wire [15:0] _T_94961; // @[Mux.scala 31:69:@39952.4]
  wire [15:0] _T_94962; // @[Mux.scala 31:69:@39953.4]
  wire [15:0] _T_94963; // @[Mux.scala 31:69:@39954.4]
  wire [15:0] _T_94964; // @[Mux.scala 31:69:@39955.4]
  wire [15:0] _T_94965; // @[Mux.scala 31:69:@39956.4]
  wire [15:0] _T_94966; // @[Mux.scala 31:69:@39957.4]
  wire [15:0] _T_94967; // @[Mux.scala 31:69:@39958.4]
  wire [15:0] _T_94968; // @[Mux.scala 31:69:@39959.4]
  wire [15:0] _T_94969; // @[Mux.scala 31:69:@39960.4]
  wire [15:0] _T_94970; // @[Mux.scala 31:69:@39961.4]
  wire [15:0] _T_94971; // @[Mux.scala 31:69:@39962.4]
  wire  _T_94972; // @[OneHot.scala 66:30:@39963.4]
  wire  _T_94973; // @[OneHot.scala 66:30:@39964.4]
  wire  _T_94974; // @[OneHot.scala 66:30:@39965.4]
  wire  _T_94975; // @[OneHot.scala 66:30:@39966.4]
  wire  _T_94976; // @[OneHot.scala 66:30:@39967.4]
  wire  _T_94977; // @[OneHot.scala 66:30:@39968.4]
  wire  _T_94978; // @[OneHot.scala 66:30:@39969.4]
  wire  _T_94979; // @[OneHot.scala 66:30:@39970.4]
  wire  _T_94980; // @[OneHot.scala 66:30:@39971.4]
  wire  _T_94981; // @[OneHot.scala 66:30:@39972.4]
  wire  _T_94982; // @[OneHot.scala 66:30:@39973.4]
  wire  _T_94983; // @[OneHot.scala 66:30:@39974.4]
  wire  _T_94984; // @[OneHot.scala 66:30:@39975.4]
  wire  _T_94985; // @[OneHot.scala 66:30:@39976.4]
  wire  _T_94986; // @[OneHot.scala 66:30:@39977.4]
  wire  _T_94987; // @[OneHot.scala 66:30:@39978.4]
  wire [15:0] _T_95028; // @[Mux.scala 31:69:@39996.4]
  wire [15:0] _T_95029; // @[Mux.scala 31:69:@39997.4]
  wire [15:0] _T_95030; // @[Mux.scala 31:69:@39998.4]
  wire [15:0] _T_95031; // @[Mux.scala 31:69:@39999.4]
  wire [15:0] _T_95032; // @[Mux.scala 31:69:@40000.4]
  wire [15:0] _T_95033; // @[Mux.scala 31:69:@40001.4]
  wire [15:0] _T_95034; // @[Mux.scala 31:69:@40002.4]
  wire [15:0] _T_95035; // @[Mux.scala 31:69:@40003.4]
  wire [15:0] _T_95036; // @[Mux.scala 31:69:@40004.4]
  wire [15:0] _T_95037; // @[Mux.scala 31:69:@40005.4]
  wire [15:0] _T_95038; // @[Mux.scala 31:69:@40006.4]
  wire [15:0] _T_95039; // @[Mux.scala 31:69:@40007.4]
  wire [15:0] _T_95040; // @[Mux.scala 31:69:@40008.4]
  wire [15:0] _T_95041; // @[Mux.scala 31:69:@40009.4]
  wire [15:0] _T_95042; // @[Mux.scala 31:69:@40010.4]
  wire [15:0] _T_95043; // @[Mux.scala 31:69:@40011.4]
  wire  _T_95044; // @[OneHot.scala 66:30:@40012.4]
  wire  _T_95045; // @[OneHot.scala 66:30:@40013.4]
  wire  _T_95046; // @[OneHot.scala 66:30:@40014.4]
  wire  _T_95047; // @[OneHot.scala 66:30:@40015.4]
  wire  _T_95048; // @[OneHot.scala 66:30:@40016.4]
  wire  _T_95049; // @[OneHot.scala 66:30:@40017.4]
  wire  _T_95050; // @[OneHot.scala 66:30:@40018.4]
  wire  _T_95051; // @[OneHot.scala 66:30:@40019.4]
  wire  _T_95052; // @[OneHot.scala 66:30:@40020.4]
  wire  _T_95053; // @[OneHot.scala 66:30:@40021.4]
  wire  _T_95054; // @[OneHot.scala 66:30:@40022.4]
  wire  _T_95055; // @[OneHot.scala 66:30:@40023.4]
  wire  _T_95056; // @[OneHot.scala 66:30:@40024.4]
  wire  _T_95057; // @[OneHot.scala 66:30:@40025.4]
  wire  _T_95058; // @[OneHot.scala 66:30:@40026.4]
  wire  _T_95059; // @[OneHot.scala 66:30:@40027.4]
  wire [15:0] _T_95100; // @[Mux.scala 31:69:@40045.4]
  wire [15:0] _T_95101; // @[Mux.scala 31:69:@40046.4]
  wire [15:0] _T_95102; // @[Mux.scala 31:69:@40047.4]
  wire [15:0] _T_95103; // @[Mux.scala 31:69:@40048.4]
  wire [15:0] _T_95104; // @[Mux.scala 31:69:@40049.4]
  wire [15:0] _T_95105; // @[Mux.scala 31:69:@40050.4]
  wire [15:0] _T_95106; // @[Mux.scala 31:69:@40051.4]
  wire [15:0] _T_95107; // @[Mux.scala 31:69:@40052.4]
  wire [15:0] _T_95108; // @[Mux.scala 31:69:@40053.4]
  wire [15:0] _T_95109; // @[Mux.scala 31:69:@40054.4]
  wire [15:0] _T_95110; // @[Mux.scala 31:69:@40055.4]
  wire [15:0] _T_95111; // @[Mux.scala 31:69:@40056.4]
  wire [15:0] _T_95112; // @[Mux.scala 31:69:@40057.4]
  wire [15:0] _T_95113; // @[Mux.scala 31:69:@40058.4]
  wire [15:0] _T_95114; // @[Mux.scala 31:69:@40059.4]
  wire [15:0] _T_95115; // @[Mux.scala 31:69:@40060.4]
  wire  _T_95116; // @[OneHot.scala 66:30:@40061.4]
  wire  _T_95117; // @[OneHot.scala 66:30:@40062.4]
  wire  _T_95118; // @[OneHot.scala 66:30:@40063.4]
  wire  _T_95119; // @[OneHot.scala 66:30:@40064.4]
  wire  _T_95120; // @[OneHot.scala 66:30:@40065.4]
  wire  _T_95121; // @[OneHot.scala 66:30:@40066.4]
  wire  _T_95122; // @[OneHot.scala 66:30:@40067.4]
  wire  _T_95123; // @[OneHot.scala 66:30:@40068.4]
  wire  _T_95124; // @[OneHot.scala 66:30:@40069.4]
  wire  _T_95125; // @[OneHot.scala 66:30:@40070.4]
  wire  _T_95126; // @[OneHot.scala 66:30:@40071.4]
  wire  _T_95127; // @[OneHot.scala 66:30:@40072.4]
  wire  _T_95128; // @[OneHot.scala 66:30:@40073.4]
  wire  _T_95129; // @[OneHot.scala 66:30:@40074.4]
  wire  _T_95130; // @[OneHot.scala 66:30:@40075.4]
  wire  _T_95131; // @[OneHot.scala 66:30:@40076.4]
  wire [15:0] _T_95172; // @[Mux.scala 31:69:@40094.4]
  wire [15:0] _T_95173; // @[Mux.scala 31:69:@40095.4]
  wire [15:0] _T_95174; // @[Mux.scala 31:69:@40096.4]
  wire [15:0] _T_95175; // @[Mux.scala 31:69:@40097.4]
  wire [15:0] _T_95176; // @[Mux.scala 31:69:@40098.4]
  wire [15:0] _T_95177; // @[Mux.scala 31:69:@40099.4]
  wire [15:0] _T_95178; // @[Mux.scala 31:69:@40100.4]
  wire [15:0] _T_95179; // @[Mux.scala 31:69:@40101.4]
  wire [15:0] _T_95180; // @[Mux.scala 31:69:@40102.4]
  wire [15:0] _T_95181; // @[Mux.scala 31:69:@40103.4]
  wire [15:0] _T_95182; // @[Mux.scala 31:69:@40104.4]
  wire [15:0] _T_95183; // @[Mux.scala 31:69:@40105.4]
  wire [15:0] _T_95184; // @[Mux.scala 31:69:@40106.4]
  wire [15:0] _T_95185; // @[Mux.scala 31:69:@40107.4]
  wire [15:0] _T_95186; // @[Mux.scala 31:69:@40108.4]
  wire [15:0] _T_95187; // @[Mux.scala 31:69:@40109.4]
  wire  _T_95188; // @[OneHot.scala 66:30:@40110.4]
  wire  _T_95189; // @[OneHot.scala 66:30:@40111.4]
  wire  _T_95190; // @[OneHot.scala 66:30:@40112.4]
  wire  _T_95191; // @[OneHot.scala 66:30:@40113.4]
  wire  _T_95192; // @[OneHot.scala 66:30:@40114.4]
  wire  _T_95193; // @[OneHot.scala 66:30:@40115.4]
  wire  _T_95194; // @[OneHot.scala 66:30:@40116.4]
  wire  _T_95195; // @[OneHot.scala 66:30:@40117.4]
  wire  _T_95196; // @[OneHot.scala 66:30:@40118.4]
  wire  _T_95197; // @[OneHot.scala 66:30:@40119.4]
  wire  _T_95198; // @[OneHot.scala 66:30:@40120.4]
  wire  _T_95199; // @[OneHot.scala 66:30:@40121.4]
  wire  _T_95200; // @[OneHot.scala 66:30:@40122.4]
  wire  _T_95201; // @[OneHot.scala 66:30:@40123.4]
  wire  _T_95202; // @[OneHot.scala 66:30:@40124.4]
  wire  _T_95203; // @[OneHot.scala 66:30:@40125.4]
  wire [15:0] _T_95244; // @[Mux.scala 31:69:@40143.4]
  wire [15:0] _T_95245; // @[Mux.scala 31:69:@40144.4]
  wire [15:0] _T_95246; // @[Mux.scala 31:69:@40145.4]
  wire [15:0] _T_95247; // @[Mux.scala 31:69:@40146.4]
  wire [15:0] _T_95248; // @[Mux.scala 31:69:@40147.4]
  wire [15:0] _T_95249; // @[Mux.scala 31:69:@40148.4]
  wire [15:0] _T_95250; // @[Mux.scala 31:69:@40149.4]
  wire [15:0] _T_95251; // @[Mux.scala 31:69:@40150.4]
  wire [15:0] _T_95252; // @[Mux.scala 31:69:@40151.4]
  wire [15:0] _T_95253; // @[Mux.scala 31:69:@40152.4]
  wire [15:0] _T_95254; // @[Mux.scala 31:69:@40153.4]
  wire [15:0] _T_95255; // @[Mux.scala 31:69:@40154.4]
  wire [15:0] _T_95256; // @[Mux.scala 31:69:@40155.4]
  wire [15:0] _T_95257; // @[Mux.scala 31:69:@40156.4]
  wire [15:0] _T_95258; // @[Mux.scala 31:69:@40157.4]
  wire [15:0] _T_95259; // @[Mux.scala 31:69:@40158.4]
  wire  _T_95260; // @[OneHot.scala 66:30:@40159.4]
  wire  _T_95261; // @[OneHot.scala 66:30:@40160.4]
  wire  _T_95262; // @[OneHot.scala 66:30:@40161.4]
  wire  _T_95263; // @[OneHot.scala 66:30:@40162.4]
  wire  _T_95264; // @[OneHot.scala 66:30:@40163.4]
  wire  _T_95265; // @[OneHot.scala 66:30:@40164.4]
  wire  _T_95266; // @[OneHot.scala 66:30:@40165.4]
  wire  _T_95267; // @[OneHot.scala 66:30:@40166.4]
  wire  _T_95268; // @[OneHot.scala 66:30:@40167.4]
  wire  _T_95269; // @[OneHot.scala 66:30:@40168.4]
  wire  _T_95270; // @[OneHot.scala 66:30:@40169.4]
  wire  _T_95271; // @[OneHot.scala 66:30:@40170.4]
  wire  _T_95272; // @[OneHot.scala 66:30:@40171.4]
  wire  _T_95273; // @[OneHot.scala 66:30:@40172.4]
  wire  _T_95274; // @[OneHot.scala 66:30:@40173.4]
  wire  _T_95275; // @[OneHot.scala 66:30:@40174.4]
  wire [15:0] _T_95316; // @[Mux.scala 31:69:@40192.4]
  wire [15:0] _T_95317; // @[Mux.scala 31:69:@40193.4]
  wire [15:0] _T_95318; // @[Mux.scala 31:69:@40194.4]
  wire [15:0] _T_95319; // @[Mux.scala 31:69:@40195.4]
  wire [15:0] _T_95320; // @[Mux.scala 31:69:@40196.4]
  wire [15:0] _T_95321; // @[Mux.scala 31:69:@40197.4]
  wire [15:0] _T_95322; // @[Mux.scala 31:69:@40198.4]
  wire [15:0] _T_95323; // @[Mux.scala 31:69:@40199.4]
  wire [15:0] _T_95324; // @[Mux.scala 31:69:@40200.4]
  wire [15:0] _T_95325; // @[Mux.scala 31:69:@40201.4]
  wire [15:0] _T_95326; // @[Mux.scala 31:69:@40202.4]
  wire [15:0] _T_95327; // @[Mux.scala 31:69:@40203.4]
  wire [15:0] _T_95328; // @[Mux.scala 31:69:@40204.4]
  wire [15:0] _T_95329; // @[Mux.scala 31:69:@40205.4]
  wire [15:0] _T_95330; // @[Mux.scala 31:69:@40206.4]
  wire [15:0] _T_95331; // @[Mux.scala 31:69:@40207.4]
  wire  _T_95332; // @[OneHot.scala 66:30:@40208.4]
  wire  _T_95333; // @[OneHot.scala 66:30:@40209.4]
  wire  _T_95334; // @[OneHot.scala 66:30:@40210.4]
  wire  _T_95335; // @[OneHot.scala 66:30:@40211.4]
  wire  _T_95336; // @[OneHot.scala 66:30:@40212.4]
  wire  _T_95337; // @[OneHot.scala 66:30:@40213.4]
  wire  _T_95338; // @[OneHot.scala 66:30:@40214.4]
  wire  _T_95339; // @[OneHot.scala 66:30:@40215.4]
  wire  _T_95340; // @[OneHot.scala 66:30:@40216.4]
  wire  _T_95341; // @[OneHot.scala 66:30:@40217.4]
  wire  _T_95342; // @[OneHot.scala 66:30:@40218.4]
  wire  _T_95343; // @[OneHot.scala 66:30:@40219.4]
  wire  _T_95344; // @[OneHot.scala 66:30:@40220.4]
  wire  _T_95345; // @[OneHot.scala 66:30:@40221.4]
  wire  _T_95346; // @[OneHot.scala 66:30:@40222.4]
  wire  _T_95347; // @[OneHot.scala 66:30:@40223.4]
  wire [15:0] _T_95388; // @[Mux.scala 31:69:@40241.4]
  wire [15:0] _T_95389; // @[Mux.scala 31:69:@40242.4]
  wire [15:0] _T_95390; // @[Mux.scala 31:69:@40243.4]
  wire [15:0] _T_95391; // @[Mux.scala 31:69:@40244.4]
  wire [15:0] _T_95392; // @[Mux.scala 31:69:@40245.4]
  wire [15:0] _T_95393; // @[Mux.scala 31:69:@40246.4]
  wire [15:0] _T_95394; // @[Mux.scala 31:69:@40247.4]
  wire [15:0] _T_95395; // @[Mux.scala 31:69:@40248.4]
  wire [15:0] _T_95396; // @[Mux.scala 31:69:@40249.4]
  wire [15:0] _T_95397; // @[Mux.scala 31:69:@40250.4]
  wire [15:0] _T_95398; // @[Mux.scala 31:69:@40251.4]
  wire [15:0] _T_95399; // @[Mux.scala 31:69:@40252.4]
  wire [15:0] _T_95400; // @[Mux.scala 31:69:@40253.4]
  wire [15:0] _T_95401; // @[Mux.scala 31:69:@40254.4]
  wire [15:0] _T_95402; // @[Mux.scala 31:69:@40255.4]
  wire [15:0] _T_95403; // @[Mux.scala 31:69:@40256.4]
  wire  _T_95404; // @[OneHot.scala 66:30:@40257.4]
  wire  _T_95405; // @[OneHot.scala 66:30:@40258.4]
  wire  _T_95406; // @[OneHot.scala 66:30:@40259.4]
  wire  _T_95407; // @[OneHot.scala 66:30:@40260.4]
  wire  _T_95408; // @[OneHot.scala 66:30:@40261.4]
  wire  _T_95409; // @[OneHot.scala 66:30:@40262.4]
  wire  _T_95410; // @[OneHot.scala 66:30:@40263.4]
  wire  _T_95411; // @[OneHot.scala 66:30:@40264.4]
  wire  _T_95412; // @[OneHot.scala 66:30:@40265.4]
  wire  _T_95413; // @[OneHot.scala 66:30:@40266.4]
  wire  _T_95414; // @[OneHot.scala 66:30:@40267.4]
  wire  _T_95415; // @[OneHot.scala 66:30:@40268.4]
  wire  _T_95416; // @[OneHot.scala 66:30:@40269.4]
  wire  _T_95417; // @[OneHot.scala 66:30:@40270.4]
  wire  _T_95418; // @[OneHot.scala 66:30:@40271.4]
  wire  _T_95419; // @[OneHot.scala 66:30:@40272.4]
  wire [7:0] _T_95484; // @[Mux.scala 19:72:@40296.4]
  wire [15:0] _T_95492; // @[Mux.scala 19:72:@40304.4]
  wire [15:0] _T_95494; // @[Mux.scala 19:72:@40305.4]
  wire [7:0] _T_95501; // @[Mux.scala 19:72:@40312.4]
  wire [15:0] _T_95509; // @[Mux.scala 19:72:@40320.4]
  wire [15:0] _T_95511; // @[Mux.scala 19:72:@40321.4]
  wire [7:0] _T_95518; // @[Mux.scala 19:72:@40328.4]
  wire [15:0] _T_95526; // @[Mux.scala 19:72:@40336.4]
  wire [15:0] _T_95528; // @[Mux.scala 19:72:@40337.4]
  wire [7:0] _T_95535; // @[Mux.scala 19:72:@40344.4]
  wire [15:0] _T_95543; // @[Mux.scala 19:72:@40352.4]
  wire [15:0] _T_95545; // @[Mux.scala 19:72:@40353.4]
  wire [7:0] _T_95552; // @[Mux.scala 19:72:@40360.4]
  wire [15:0] _T_95560; // @[Mux.scala 19:72:@40368.4]
  wire [15:0] _T_95562; // @[Mux.scala 19:72:@40369.4]
  wire [7:0] _T_95569; // @[Mux.scala 19:72:@40376.4]
  wire [15:0] _T_95577; // @[Mux.scala 19:72:@40384.4]
  wire [15:0] _T_95579; // @[Mux.scala 19:72:@40385.4]
  wire [7:0] _T_95586; // @[Mux.scala 19:72:@40392.4]
  wire [15:0] _T_95594; // @[Mux.scala 19:72:@40400.4]
  wire [15:0] _T_95596; // @[Mux.scala 19:72:@40401.4]
  wire [7:0] _T_95603; // @[Mux.scala 19:72:@40408.4]
  wire [15:0] _T_95611; // @[Mux.scala 19:72:@40416.4]
  wire [15:0] _T_95613; // @[Mux.scala 19:72:@40417.4]
  wire [7:0] _T_95620; // @[Mux.scala 19:72:@40424.4]
  wire [15:0] _T_95628; // @[Mux.scala 19:72:@40432.4]
  wire [15:0] _T_95630; // @[Mux.scala 19:72:@40433.4]
  wire [7:0] _T_95637; // @[Mux.scala 19:72:@40440.4]
  wire [15:0] _T_95645; // @[Mux.scala 19:72:@40448.4]
  wire [15:0] _T_95647; // @[Mux.scala 19:72:@40449.4]
  wire [7:0] _T_95654; // @[Mux.scala 19:72:@40456.4]
  wire [15:0] _T_95662; // @[Mux.scala 19:72:@40464.4]
  wire [15:0] _T_95664; // @[Mux.scala 19:72:@40465.4]
  wire [7:0] _T_95671; // @[Mux.scala 19:72:@40472.4]
  wire [15:0] _T_95679; // @[Mux.scala 19:72:@40480.4]
  wire [15:0] _T_95681; // @[Mux.scala 19:72:@40481.4]
  wire [7:0] _T_95688; // @[Mux.scala 19:72:@40488.4]
  wire [15:0] _T_95696; // @[Mux.scala 19:72:@40496.4]
  wire [15:0] _T_95698; // @[Mux.scala 19:72:@40497.4]
  wire [7:0] _T_95705; // @[Mux.scala 19:72:@40504.4]
  wire [15:0] _T_95713; // @[Mux.scala 19:72:@40512.4]
  wire [15:0] _T_95715; // @[Mux.scala 19:72:@40513.4]
  wire [7:0] _T_95722; // @[Mux.scala 19:72:@40520.4]
  wire [15:0] _T_95730; // @[Mux.scala 19:72:@40528.4]
  wire [15:0] _T_95732; // @[Mux.scala 19:72:@40529.4]
  wire [7:0] _T_95739; // @[Mux.scala 19:72:@40536.4]
  wire [15:0] _T_95747; // @[Mux.scala 19:72:@40544.4]
  wire [15:0] _T_95749; // @[Mux.scala 19:72:@40545.4]
  wire [15:0] _T_95750; // @[Mux.scala 19:72:@40546.4]
  wire [15:0] _T_95751; // @[Mux.scala 19:72:@40547.4]
  wire [15:0] _T_95752; // @[Mux.scala 19:72:@40548.4]
  wire [15:0] _T_95753; // @[Mux.scala 19:72:@40549.4]
  wire [15:0] _T_95754; // @[Mux.scala 19:72:@40550.4]
  wire [15:0] _T_95755; // @[Mux.scala 19:72:@40551.4]
  wire [15:0] _T_95756; // @[Mux.scala 19:72:@40552.4]
  wire [15:0] _T_95757; // @[Mux.scala 19:72:@40553.4]
  wire [15:0] _T_95758; // @[Mux.scala 19:72:@40554.4]
  wire [15:0] _T_95759; // @[Mux.scala 19:72:@40555.4]
  wire [15:0] _T_95760; // @[Mux.scala 19:72:@40556.4]
  wire [15:0] _T_95761; // @[Mux.scala 19:72:@40557.4]
  wire [15:0] _T_95762; // @[Mux.scala 19:72:@40558.4]
  wire [15:0] _T_95763; // @[Mux.scala 19:72:@40559.4]
  wire [15:0] _T_95764; // @[Mux.scala 19:72:@40560.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@40564.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@40566.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@40568.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@40570.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@40572.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@40574.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@40576.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@40578.4]
  wire  inputPriorityPorts_0_8; // @[Mux.scala 19:72:@40580.4]
  wire  inputPriorityPorts_0_9; // @[Mux.scala 19:72:@40582.4]
  wire  inputPriorityPorts_0_10; // @[Mux.scala 19:72:@40584.4]
  wire  inputPriorityPorts_0_11; // @[Mux.scala 19:72:@40586.4]
  wire  inputPriorityPorts_0_12; // @[Mux.scala 19:72:@40588.4]
  wire  inputPriorityPorts_0_13; // @[Mux.scala 19:72:@40590.4]
  wire  inputPriorityPorts_0_14; // @[Mux.scala 19:72:@40592.4]
  wire  inputPriorityPorts_0_15; // @[Mux.scala 19:72:@40594.4]
  wire [15:0] _T_95966; // @[Mux.scala 31:69:@40648.4]
  wire [15:0] _T_95967; // @[Mux.scala 31:69:@40649.4]
  wire [15:0] _T_95968; // @[Mux.scala 31:69:@40650.4]
  wire [15:0] _T_95969; // @[Mux.scala 31:69:@40651.4]
  wire [15:0] _T_95970; // @[Mux.scala 31:69:@40652.4]
  wire [15:0] _T_95971; // @[Mux.scala 31:69:@40653.4]
  wire [15:0] _T_95972; // @[Mux.scala 31:69:@40654.4]
  wire [15:0] _T_95973; // @[Mux.scala 31:69:@40655.4]
  wire [15:0] _T_95974; // @[Mux.scala 31:69:@40656.4]
  wire [15:0] _T_95975; // @[Mux.scala 31:69:@40657.4]
  wire [15:0] _T_95976; // @[Mux.scala 31:69:@40658.4]
  wire [15:0] _T_95977; // @[Mux.scala 31:69:@40659.4]
  wire [15:0] _T_95978; // @[Mux.scala 31:69:@40660.4]
  wire [15:0] _T_95979; // @[Mux.scala 31:69:@40661.4]
  wire [15:0] _T_95980; // @[Mux.scala 31:69:@40662.4]
  wire [15:0] _T_95981; // @[Mux.scala 31:69:@40663.4]
  wire  _T_95982; // @[OneHot.scala 66:30:@40664.4]
  wire  _T_95983; // @[OneHot.scala 66:30:@40665.4]
  wire  _T_95984; // @[OneHot.scala 66:30:@40666.4]
  wire  _T_95985; // @[OneHot.scala 66:30:@40667.4]
  wire  _T_95986; // @[OneHot.scala 66:30:@40668.4]
  wire  _T_95987; // @[OneHot.scala 66:30:@40669.4]
  wire  _T_95988; // @[OneHot.scala 66:30:@40670.4]
  wire  _T_95989; // @[OneHot.scala 66:30:@40671.4]
  wire  _T_95990; // @[OneHot.scala 66:30:@40672.4]
  wire  _T_95991; // @[OneHot.scala 66:30:@40673.4]
  wire  _T_95992; // @[OneHot.scala 66:30:@40674.4]
  wire  _T_95993; // @[OneHot.scala 66:30:@40675.4]
  wire  _T_95994; // @[OneHot.scala 66:30:@40676.4]
  wire  _T_95995; // @[OneHot.scala 66:30:@40677.4]
  wire  _T_95996; // @[OneHot.scala 66:30:@40678.4]
  wire  _T_95997; // @[OneHot.scala 66:30:@40679.4]
  wire [15:0] _T_96038; // @[Mux.scala 31:69:@40697.4]
  wire [15:0] _T_96039; // @[Mux.scala 31:69:@40698.4]
  wire [15:0] _T_96040; // @[Mux.scala 31:69:@40699.4]
  wire [15:0] _T_96041; // @[Mux.scala 31:69:@40700.4]
  wire [15:0] _T_96042; // @[Mux.scala 31:69:@40701.4]
  wire [15:0] _T_96043; // @[Mux.scala 31:69:@40702.4]
  wire [15:0] _T_96044; // @[Mux.scala 31:69:@40703.4]
  wire [15:0] _T_96045; // @[Mux.scala 31:69:@40704.4]
  wire [15:0] _T_96046; // @[Mux.scala 31:69:@40705.4]
  wire [15:0] _T_96047; // @[Mux.scala 31:69:@40706.4]
  wire [15:0] _T_96048; // @[Mux.scala 31:69:@40707.4]
  wire [15:0] _T_96049; // @[Mux.scala 31:69:@40708.4]
  wire [15:0] _T_96050; // @[Mux.scala 31:69:@40709.4]
  wire [15:0] _T_96051; // @[Mux.scala 31:69:@40710.4]
  wire [15:0] _T_96052; // @[Mux.scala 31:69:@40711.4]
  wire [15:0] _T_96053; // @[Mux.scala 31:69:@40712.4]
  wire  _T_96054; // @[OneHot.scala 66:30:@40713.4]
  wire  _T_96055; // @[OneHot.scala 66:30:@40714.4]
  wire  _T_96056; // @[OneHot.scala 66:30:@40715.4]
  wire  _T_96057; // @[OneHot.scala 66:30:@40716.4]
  wire  _T_96058; // @[OneHot.scala 66:30:@40717.4]
  wire  _T_96059; // @[OneHot.scala 66:30:@40718.4]
  wire  _T_96060; // @[OneHot.scala 66:30:@40719.4]
  wire  _T_96061; // @[OneHot.scala 66:30:@40720.4]
  wire  _T_96062; // @[OneHot.scala 66:30:@40721.4]
  wire  _T_96063; // @[OneHot.scala 66:30:@40722.4]
  wire  _T_96064; // @[OneHot.scala 66:30:@40723.4]
  wire  _T_96065; // @[OneHot.scala 66:30:@40724.4]
  wire  _T_96066; // @[OneHot.scala 66:30:@40725.4]
  wire  _T_96067; // @[OneHot.scala 66:30:@40726.4]
  wire  _T_96068; // @[OneHot.scala 66:30:@40727.4]
  wire  _T_96069; // @[OneHot.scala 66:30:@40728.4]
  wire [15:0] _T_96110; // @[Mux.scala 31:69:@40746.4]
  wire [15:0] _T_96111; // @[Mux.scala 31:69:@40747.4]
  wire [15:0] _T_96112; // @[Mux.scala 31:69:@40748.4]
  wire [15:0] _T_96113; // @[Mux.scala 31:69:@40749.4]
  wire [15:0] _T_96114; // @[Mux.scala 31:69:@40750.4]
  wire [15:0] _T_96115; // @[Mux.scala 31:69:@40751.4]
  wire [15:0] _T_96116; // @[Mux.scala 31:69:@40752.4]
  wire [15:0] _T_96117; // @[Mux.scala 31:69:@40753.4]
  wire [15:0] _T_96118; // @[Mux.scala 31:69:@40754.4]
  wire [15:0] _T_96119; // @[Mux.scala 31:69:@40755.4]
  wire [15:0] _T_96120; // @[Mux.scala 31:69:@40756.4]
  wire [15:0] _T_96121; // @[Mux.scala 31:69:@40757.4]
  wire [15:0] _T_96122; // @[Mux.scala 31:69:@40758.4]
  wire [15:0] _T_96123; // @[Mux.scala 31:69:@40759.4]
  wire [15:0] _T_96124; // @[Mux.scala 31:69:@40760.4]
  wire [15:0] _T_96125; // @[Mux.scala 31:69:@40761.4]
  wire  _T_96126; // @[OneHot.scala 66:30:@40762.4]
  wire  _T_96127; // @[OneHot.scala 66:30:@40763.4]
  wire  _T_96128; // @[OneHot.scala 66:30:@40764.4]
  wire  _T_96129; // @[OneHot.scala 66:30:@40765.4]
  wire  _T_96130; // @[OneHot.scala 66:30:@40766.4]
  wire  _T_96131; // @[OneHot.scala 66:30:@40767.4]
  wire  _T_96132; // @[OneHot.scala 66:30:@40768.4]
  wire  _T_96133; // @[OneHot.scala 66:30:@40769.4]
  wire  _T_96134; // @[OneHot.scala 66:30:@40770.4]
  wire  _T_96135; // @[OneHot.scala 66:30:@40771.4]
  wire  _T_96136; // @[OneHot.scala 66:30:@40772.4]
  wire  _T_96137; // @[OneHot.scala 66:30:@40773.4]
  wire  _T_96138; // @[OneHot.scala 66:30:@40774.4]
  wire  _T_96139; // @[OneHot.scala 66:30:@40775.4]
  wire  _T_96140; // @[OneHot.scala 66:30:@40776.4]
  wire  _T_96141; // @[OneHot.scala 66:30:@40777.4]
  wire [15:0] _T_96182; // @[Mux.scala 31:69:@40795.4]
  wire [15:0] _T_96183; // @[Mux.scala 31:69:@40796.4]
  wire [15:0] _T_96184; // @[Mux.scala 31:69:@40797.4]
  wire [15:0] _T_96185; // @[Mux.scala 31:69:@40798.4]
  wire [15:0] _T_96186; // @[Mux.scala 31:69:@40799.4]
  wire [15:0] _T_96187; // @[Mux.scala 31:69:@40800.4]
  wire [15:0] _T_96188; // @[Mux.scala 31:69:@40801.4]
  wire [15:0] _T_96189; // @[Mux.scala 31:69:@40802.4]
  wire [15:0] _T_96190; // @[Mux.scala 31:69:@40803.4]
  wire [15:0] _T_96191; // @[Mux.scala 31:69:@40804.4]
  wire [15:0] _T_96192; // @[Mux.scala 31:69:@40805.4]
  wire [15:0] _T_96193; // @[Mux.scala 31:69:@40806.4]
  wire [15:0] _T_96194; // @[Mux.scala 31:69:@40807.4]
  wire [15:0] _T_96195; // @[Mux.scala 31:69:@40808.4]
  wire [15:0] _T_96196; // @[Mux.scala 31:69:@40809.4]
  wire [15:0] _T_96197; // @[Mux.scala 31:69:@40810.4]
  wire  _T_96198; // @[OneHot.scala 66:30:@40811.4]
  wire  _T_96199; // @[OneHot.scala 66:30:@40812.4]
  wire  _T_96200; // @[OneHot.scala 66:30:@40813.4]
  wire  _T_96201; // @[OneHot.scala 66:30:@40814.4]
  wire  _T_96202; // @[OneHot.scala 66:30:@40815.4]
  wire  _T_96203; // @[OneHot.scala 66:30:@40816.4]
  wire  _T_96204; // @[OneHot.scala 66:30:@40817.4]
  wire  _T_96205; // @[OneHot.scala 66:30:@40818.4]
  wire  _T_96206; // @[OneHot.scala 66:30:@40819.4]
  wire  _T_96207; // @[OneHot.scala 66:30:@40820.4]
  wire  _T_96208; // @[OneHot.scala 66:30:@40821.4]
  wire  _T_96209; // @[OneHot.scala 66:30:@40822.4]
  wire  _T_96210; // @[OneHot.scala 66:30:@40823.4]
  wire  _T_96211; // @[OneHot.scala 66:30:@40824.4]
  wire  _T_96212; // @[OneHot.scala 66:30:@40825.4]
  wire  _T_96213; // @[OneHot.scala 66:30:@40826.4]
  wire [15:0] _T_96254; // @[Mux.scala 31:69:@40844.4]
  wire [15:0] _T_96255; // @[Mux.scala 31:69:@40845.4]
  wire [15:0] _T_96256; // @[Mux.scala 31:69:@40846.4]
  wire [15:0] _T_96257; // @[Mux.scala 31:69:@40847.4]
  wire [15:0] _T_96258; // @[Mux.scala 31:69:@40848.4]
  wire [15:0] _T_96259; // @[Mux.scala 31:69:@40849.4]
  wire [15:0] _T_96260; // @[Mux.scala 31:69:@40850.4]
  wire [15:0] _T_96261; // @[Mux.scala 31:69:@40851.4]
  wire [15:0] _T_96262; // @[Mux.scala 31:69:@40852.4]
  wire [15:0] _T_96263; // @[Mux.scala 31:69:@40853.4]
  wire [15:0] _T_96264; // @[Mux.scala 31:69:@40854.4]
  wire [15:0] _T_96265; // @[Mux.scala 31:69:@40855.4]
  wire [15:0] _T_96266; // @[Mux.scala 31:69:@40856.4]
  wire [15:0] _T_96267; // @[Mux.scala 31:69:@40857.4]
  wire [15:0] _T_96268; // @[Mux.scala 31:69:@40858.4]
  wire [15:0] _T_96269; // @[Mux.scala 31:69:@40859.4]
  wire  _T_96270; // @[OneHot.scala 66:30:@40860.4]
  wire  _T_96271; // @[OneHot.scala 66:30:@40861.4]
  wire  _T_96272; // @[OneHot.scala 66:30:@40862.4]
  wire  _T_96273; // @[OneHot.scala 66:30:@40863.4]
  wire  _T_96274; // @[OneHot.scala 66:30:@40864.4]
  wire  _T_96275; // @[OneHot.scala 66:30:@40865.4]
  wire  _T_96276; // @[OneHot.scala 66:30:@40866.4]
  wire  _T_96277; // @[OneHot.scala 66:30:@40867.4]
  wire  _T_96278; // @[OneHot.scala 66:30:@40868.4]
  wire  _T_96279; // @[OneHot.scala 66:30:@40869.4]
  wire  _T_96280; // @[OneHot.scala 66:30:@40870.4]
  wire  _T_96281; // @[OneHot.scala 66:30:@40871.4]
  wire  _T_96282; // @[OneHot.scala 66:30:@40872.4]
  wire  _T_96283; // @[OneHot.scala 66:30:@40873.4]
  wire  _T_96284; // @[OneHot.scala 66:30:@40874.4]
  wire  _T_96285; // @[OneHot.scala 66:30:@40875.4]
  wire [15:0] _T_96326; // @[Mux.scala 31:69:@40893.4]
  wire [15:0] _T_96327; // @[Mux.scala 31:69:@40894.4]
  wire [15:0] _T_96328; // @[Mux.scala 31:69:@40895.4]
  wire [15:0] _T_96329; // @[Mux.scala 31:69:@40896.4]
  wire [15:0] _T_96330; // @[Mux.scala 31:69:@40897.4]
  wire [15:0] _T_96331; // @[Mux.scala 31:69:@40898.4]
  wire [15:0] _T_96332; // @[Mux.scala 31:69:@40899.4]
  wire [15:0] _T_96333; // @[Mux.scala 31:69:@40900.4]
  wire [15:0] _T_96334; // @[Mux.scala 31:69:@40901.4]
  wire [15:0] _T_96335; // @[Mux.scala 31:69:@40902.4]
  wire [15:0] _T_96336; // @[Mux.scala 31:69:@40903.4]
  wire [15:0] _T_96337; // @[Mux.scala 31:69:@40904.4]
  wire [15:0] _T_96338; // @[Mux.scala 31:69:@40905.4]
  wire [15:0] _T_96339; // @[Mux.scala 31:69:@40906.4]
  wire [15:0] _T_96340; // @[Mux.scala 31:69:@40907.4]
  wire [15:0] _T_96341; // @[Mux.scala 31:69:@40908.4]
  wire  _T_96342; // @[OneHot.scala 66:30:@40909.4]
  wire  _T_96343; // @[OneHot.scala 66:30:@40910.4]
  wire  _T_96344; // @[OneHot.scala 66:30:@40911.4]
  wire  _T_96345; // @[OneHot.scala 66:30:@40912.4]
  wire  _T_96346; // @[OneHot.scala 66:30:@40913.4]
  wire  _T_96347; // @[OneHot.scala 66:30:@40914.4]
  wire  _T_96348; // @[OneHot.scala 66:30:@40915.4]
  wire  _T_96349; // @[OneHot.scala 66:30:@40916.4]
  wire  _T_96350; // @[OneHot.scala 66:30:@40917.4]
  wire  _T_96351; // @[OneHot.scala 66:30:@40918.4]
  wire  _T_96352; // @[OneHot.scala 66:30:@40919.4]
  wire  _T_96353; // @[OneHot.scala 66:30:@40920.4]
  wire  _T_96354; // @[OneHot.scala 66:30:@40921.4]
  wire  _T_96355; // @[OneHot.scala 66:30:@40922.4]
  wire  _T_96356; // @[OneHot.scala 66:30:@40923.4]
  wire  _T_96357; // @[OneHot.scala 66:30:@40924.4]
  wire [15:0] _T_96398; // @[Mux.scala 31:69:@40942.4]
  wire [15:0] _T_96399; // @[Mux.scala 31:69:@40943.4]
  wire [15:0] _T_96400; // @[Mux.scala 31:69:@40944.4]
  wire [15:0] _T_96401; // @[Mux.scala 31:69:@40945.4]
  wire [15:0] _T_96402; // @[Mux.scala 31:69:@40946.4]
  wire [15:0] _T_96403; // @[Mux.scala 31:69:@40947.4]
  wire [15:0] _T_96404; // @[Mux.scala 31:69:@40948.4]
  wire [15:0] _T_96405; // @[Mux.scala 31:69:@40949.4]
  wire [15:0] _T_96406; // @[Mux.scala 31:69:@40950.4]
  wire [15:0] _T_96407; // @[Mux.scala 31:69:@40951.4]
  wire [15:0] _T_96408; // @[Mux.scala 31:69:@40952.4]
  wire [15:0] _T_96409; // @[Mux.scala 31:69:@40953.4]
  wire [15:0] _T_96410; // @[Mux.scala 31:69:@40954.4]
  wire [15:0] _T_96411; // @[Mux.scala 31:69:@40955.4]
  wire [15:0] _T_96412; // @[Mux.scala 31:69:@40956.4]
  wire [15:0] _T_96413; // @[Mux.scala 31:69:@40957.4]
  wire  _T_96414; // @[OneHot.scala 66:30:@40958.4]
  wire  _T_96415; // @[OneHot.scala 66:30:@40959.4]
  wire  _T_96416; // @[OneHot.scala 66:30:@40960.4]
  wire  _T_96417; // @[OneHot.scala 66:30:@40961.4]
  wire  _T_96418; // @[OneHot.scala 66:30:@40962.4]
  wire  _T_96419; // @[OneHot.scala 66:30:@40963.4]
  wire  _T_96420; // @[OneHot.scala 66:30:@40964.4]
  wire  _T_96421; // @[OneHot.scala 66:30:@40965.4]
  wire  _T_96422; // @[OneHot.scala 66:30:@40966.4]
  wire  _T_96423; // @[OneHot.scala 66:30:@40967.4]
  wire  _T_96424; // @[OneHot.scala 66:30:@40968.4]
  wire  _T_96425; // @[OneHot.scala 66:30:@40969.4]
  wire  _T_96426; // @[OneHot.scala 66:30:@40970.4]
  wire  _T_96427; // @[OneHot.scala 66:30:@40971.4]
  wire  _T_96428; // @[OneHot.scala 66:30:@40972.4]
  wire  _T_96429; // @[OneHot.scala 66:30:@40973.4]
  wire [15:0] _T_96470; // @[Mux.scala 31:69:@40991.4]
  wire [15:0] _T_96471; // @[Mux.scala 31:69:@40992.4]
  wire [15:0] _T_96472; // @[Mux.scala 31:69:@40993.4]
  wire [15:0] _T_96473; // @[Mux.scala 31:69:@40994.4]
  wire [15:0] _T_96474; // @[Mux.scala 31:69:@40995.4]
  wire [15:0] _T_96475; // @[Mux.scala 31:69:@40996.4]
  wire [15:0] _T_96476; // @[Mux.scala 31:69:@40997.4]
  wire [15:0] _T_96477; // @[Mux.scala 31:69:@40998.4]
  wire [15:0] _T_96478; // @[Mux.scala 31:69:@40999.4]
  wire [15:0] _T_96479; // @[Mux.scala 31:69:@41000.4]
  wire [15:0] _T_96480; // @[Mux.scala 31:69:@41001.4]
  wire [15:0] _T_96481; // @[Mux.scala 31:69:@41002.4]
  wire [15:0] _T_96482; // @[Mux.scala 31:69:@41003.4]
  wire [15:0] _T_96483; // @[Mux.scala 31:69:@41004.4]
  wire [15:0] _T_96484; // @[Mux.scala 31:69:@41005.4]
  wire [15:0] _T_96485; // @[Mux.scala 31:69:@41006.4]
  wire  _T_96486; // @[OneHot.scala 66:30:@41007.4]
  wire  _T_96487; // @[OneHot.scala 66:30:@41008.4]
  wire  _T_96488; // @[OneHot.scala 66:30:@41009.4]
  wire  _T_96489; // @[OneHot.scala 66:30:@41010.4]
  wire  _T_96490; // @[OneHot.scala 66:30:@41011.4]
  wire  _T_96491; // @[OneHot.scala 66:30:@41012.4]
  wire  _T_96492; // @[OneHot.scala 66:30:@41013.4]
  wire  _T_96493; // @[OneHot.scala 66:30:@41014.4]
  wire  _T_96494; // @[OneHot.scala 66:30:@41015.4]
  wire  _T_96495; // @[OneHot.scala 66:30:@41016.4]
  wire  _T_96496; // @[OneHot.scala 66:30:@41017.4]
  wire  _T_96497; // @[OneHot.scala 66:30:@41018.4]
  wire  _T_96498; // @[OneHot.scala 66:30:@41019.4]
  wire  _T_96499; // @[OneHot.scala 66:30:@41020.4]
  wire  _T_96500; // @[OneHot.scala 66:30:@41021.4]
  wire  _T_96501; // @[OneHot.scala 66:30:@41022.4]
  wire [15:0] _T_96542; // @[Mux.scala 31:69:@41040.4]
  wire [15:0] _T_96543; // @[Mux.scala 31:69:@41041.4]
  wire [15:0] _T_96544; // @[Mux.scala 31:69:@41042.4]
  wire [15:0] _T_96545; // @[Mux.scala 31:69:@41043.4]
  wire [15:0] _T_96546; // @[Mux.scala 31:69:@41044.4]
  wire [15:0] _T_96547; // @[Mux.scala 31:69:@41045.4]
  wire [15:0] _T_96548; // @[Mux.scala 31:69:@41046.4]
  wire [15:0] _T_96549; // @[Mux.scala 31:69:@41047.4]
  wire [15:0] _T_96550; // @[Mux.scala 31:69:@41048.4]
  wire [15:0] _T_96551; // @[Mux.scala 31:69:@41049.4]
  wire [15:0] _T_96552; // @[Mux.scala 31:69:@41050.4]
  wire [15:0] _T_96553; // @[Mux.scala 31:69:@41051.4]
  wire [15:0] _T_96554; // @[Mux.scala 31:69:@41052.4]
  wire [15:0] _T_96555; // @[Mux.scala 31:69:@41053.4]
  wire [15:0] _T_96556; // @[Mux.scala 31:69:@41054.4]
  wire [15:0] _T_96557; // @[Mux.scala 31:69:@41055.4]
  wire  _T_96558; // @[OneHot.scala 66:30:@41056.4]
  wire  _T_96559; // @[OneHot.scala 66:30:@41057.4]
  wire  _T_96560; // @[OneHot.scala 66:30:@41058.4]
  wire  _T_96561; // @[OneHot.scala 66:30:@41059.4]
  wire  _T_96562; // @[OneHot.scala 66:30:@41060.4]
  wire  _T_96563; // @[OneHot.scala 66:30:@41061.4]
  wire  _T_96564; // @[OneHot.scala 66:30:@41062.4]
  wire  _T_96565; // @[OneHot.scala 66:30:@41063.4]
  wire  _T_96566; // @[OneHot.scala 66:30:@41064.4]
  wire  _T_96567; // @[OneHot.scala 66:30:@41065.4]
  wire  _T_96568; // @[OneHot.scala 66:30:@41066.4]
  wire  _T_96569; // @[OneHot.scala 66:30:@41067.4]
  wire  _T_96570; // @[OneHot.scala 66:30:@41068.4]
  wire  _T_96571; // @[OneHot.scala 66:30:@41069.4]
  wire  _T_96572; // @[OneHot.scala 66:30:@41070.4]
  wire  _T_96573; // @[OneHot.scala 66:30:@41071.4]
  wire [15:0] _T_96614; // @[Mux.scala 31:69:@41089.4]
  wire [15:0] _T_96615; // @[Mux.scala 31:69:@41090.4]
  wire [15:0] _T_96616; // @[Mux.scala 31:69:@41091.4]
  wire [15:0] _T_96617; // @[Mux.scala 31:69:@41092.4]
  wire [15:0] _T_96618; // @[Mux.scala 31:69:@41093.4]
  wire [15:0] _T_96619; // @[Mux.scala 31:69:@41094.4]
  wire [15:0] _T_96620; // @[Mux.scala 31:69:@41095.4]
  wire [15:0] _T_96621; // @[Mux.scala 31:69:@41096.4]
  wire [15:0] _T_96622; // @[Mux.scala 31:69:@41097.4]
  wire [15:0] _T_96623; // @[Mux.scala 31:69:@41098.4]
  wire [15:0] _T_96624; // @[Mux.scala 31:69:@41099.4]
  wire [15:0] _T_96625; // @[Mux.scala 31:69:@41100.4]
  wire [15:0] _T_96626; // @[Mux.scala 31:69:@41101.4]
  wire [15:0] _T_96627; // @[Mux.scala 31:69:@41102.4]
  wire [15:0] _T_96628; // @[Mux.scala 31:69:@41103.4]
  wire [15:0] _T_96629; // @[Mux.scala 31:69:@41104.4]
  wire  _T_96630; // @[OneHot.scala 66:30:@41105.4]
  wire  _T_96631; // @[OneHot.scala 66:30:@41106.4]
  wire  _T_96632; // @[OneHot.scala 66:30:@41107.4]
  wire  _T_96633; // @[OneHot.scala 66:30:@41108.4]
  wire  _T_96634; // @[OneHot.scala 66:30:@41109.4]
  wire  _T_96635; // @[OneHot.scala 66:30:@41110.4]
  wire  _T_96636; // @[OneHot.scala 66:30:@41111.4]
  wire  _T_96637; // @[OneHot.scala 66:30:@41112.4]
  wire  _T_96638; // @[OneHot.scala 66:30:@41113.4]
  wire  _T_96639; // @[OneHot.scala 66:30:@41114.4]
  wire  _T_96640; // @[OneHot.scala 66:30:@41115.4]
  wire  _T_96641; // @[OneHot.scala 66:30:@41116.4]
  wire  _T_96642; // @[OneHot.scala 66:30:@41117.4]
  wire  _T_96643; // @[OneHot.scala 66:30:@41118.4]
  wire  _T_96644; // @[OneHot.scala 66:30:@41119.4]
  wire  _T_96645; // @[OneHot.scala 66:30:@41120.4]
  wire [15:0] _T_96686; // @[Mux.scala 31:69:@41138.4]
  wire [15:0] _T_96687; // @[Mux.scala 31:69:@41139.4]
  wire [15:0] _T_96688; // @[Mux.scala 31:69:@41140.4]
  wire [15:0] _T_96689; // @[Mux.scala 31:69:@41141.4]
  wire [15:0] _T_96690; // @[Mux.scala 31:69:@41142.4]
  wire [15:0] _T_96691; // @[Mux.scala 31:69:@41143.4]
  wire [15:0] _T_96692; // @[Mux.scala 31:69:@41144.4]
  wire [15:0] _T_96693; // @[Mux.scala 31:69:@41145.4]
  wire [15:0] _T_96694; // @[Mux.scala 31:69:@41146.4]
  wire [15:0] _T_96695; // @[Mux.scala 31:69:@41147.4]
  wire [15:0] _T_96696; // @[Mux.scala 31:69:@41148.4]
  wire [15:0] _T_96697; // @[Mux.scala 31:69:@41149.4]
  wire [15:0] _T_96698; // @[Mux.scala 31:69:@41150.4]
  wire [15:0] _T_96699; // @[Mux.scala 31:69:@41151.4]
  wire [15:0] _T_96700; // @[Mux.scala 31:69:@41152.4]
  wire [15:0] _T_96701; // @[Mux.scala 31:69:@41153.4]
  wire  _T_96702; // @[OneHot.scala 66:30:@41154.4]
  wire  _T_96703; // @[OneHot.scala 66:30:@41155.4]
  wire  _T_96704; // @[OneHot.scala 66:30:@41156.4]
  wire  _T_96705; // @[OneHot.scala 66:30:@41157.4]
  wire  _T_96706; // @[OneHot.scala 66:30:@41158.4]
  wire  _T_96707; // @[OneHot.scala 66:30:@41159.4]
  wire  _T_96708; // @[OneHot.scala 66:30:@41160.4]
  wire  _T_96709; // @[OneHot.scala 66:30:@41161.4]
  wire  _T_96710; // @[OneHot.scala 66:30:@41162.4]
  wire  _T_96711; // @[OneHot.scala 66:30:@41163.4]
  wire  _T_96712; // @[OneHot.scala 66:30:@41164.4]
  wire  _T_96713; // @[OneHot.scala 66:30:@41165.4]
  wire  _T_96714; // @[OneHot.scala 66:30:@41166.4]
  wire  _T_96715; // @[OneHot.scala 66:30:@41167.4]
  wire  _T_96716; // @[OneHot.scala 66:30:@41168.4]
  wire  _T_96717; // @[OneHot.scala 66:30:@41169.4]
  wire [15:0] _T_96758; // @[Mux.scala 31:69:@41187.4]
  wire [15:0] _T_96759; // @[Mux.scala 31:69:@41188.4]
  wire [15:0] _T_96760; // @[Mux.scala 31:69:@41189.4]
  wire [15:0] _T_96761; // @[Mux.scala 31:69:@41190.4]
  wire [15:0] _T_96762; // @[Mux.scala 31:69:@41191.4]
  wire [15:0] _T_96763; // @[Mux.scala 31:69:@41192.4]
  wire [15:0] _T_96764; // @[Mux.scala 31:69:@41193.4]
  wire [15:0] _T_96765; // @[Mux.scala 31:69:@41194.4]
  wire [15:0] _T_96766; // @[Mux.scala 31:69:@41195.4]
  wire [15:0] _T_96767; // @[Mux.scala 31:69:@41196.4]
  wire [15:0] _T_96768; // @[Mux.scala 31:69:@41197.4]
  wire [15:0] _T_96769; // @[Mux.scala 31:69:@41198.4]
  wire [15:0] _T_96770; // @[Mux.scala 31:69:@41199.4]
  wire [15:0] _T_96771; // @[Mux.scala 31:69:@41200.4]
  wire [15:0] _T_96772; // @[Mux.scala 31:69:@41201.4]
  wire [15:0] _T_96773; // @[Mux.scala 31:69:@41202.4]
  wire  _T_96774; // @[OneHot.scala 66:30:@41203.4]
  wire  _T_96775; // @[OneHot.scala 66:30:@41204.4]
  wire  _T_96776; // @[OneHot.scala 66:30:@41205.4]
  wire  _T_96777; // @[OneHot.scala 66:30:@41206.4]
  wire  _T_96778; // @[OneHot.scala 66:30:@41207.4]
  wire  _T_96779; // @[OneHot.scala 66:30:@41208.4]
  wire  _T_96780; // @[OneHot.scala 66:30:@41209.4]
  wire  _T_96781; // @[OneHot.scala 66:30:@41210.4]
  wire  _T_96782; // @[OneHot.scala 66:30:@41211.4]
  wire  _T_96783; // @[OneHot.scala 66:30:@41212.4]
  wire  _T_96784; // @[OneHot.scala 66:30:@41213.4]
  wire  _T_96785; // @[OneHot.scala 66:30:@41214.4]
  wire  _T_96786; // @[OneHot.scala 66:30:@41215.4]
  wire  _T_96787; // @[OneHot.scala 66:30:@41216.4]
  wire  _T_96788; // @[OneHot.scala 66:30:@41217.4]
  wire  _T_96789; // @[OneHot.scala 66:30:@41218.4]
  wire [15:0] _T_96830; // @[Mux.scala 31:69:@41236.4]
  wire [15:0] _T_96831; // @[Mux.scala 31:69:@41237.4]
  wire [15:0] _T_96832; // @[Mux.scala 31:69:@41238.4]
  wire [15:0] _T_96833; // @[Mux.scala 31:69:@41239.4]
  wire [15:0] _T_96834; // @[Mux.scala 31:69:@41240.4]
  wire [15:0] _T_96835; // @[Mux.scala 31:69:@41241.4]
  wire [15:0] _T_96836; // @[Mux.scala 31:69:@41242.4]
  wire [15:0] _T_96837; // @[Mux.scala 31:69:@41243.4]
  wire [15:0] _T_96838; // @[Mux.scala 31:69:@41244.4]
  wire [15:0] _T_96839; // @[Mux.scala 31:69:@41245.4]
  wire [15:0] _T_96840; // @[Mux.scala 31:69:@41246.4]
  wire [15:0] _T_96841; // @[Mux.scala 31:69:@41247.4]
  wire [15:0] _T_96842; // @[Mux.scala 31:69:@41248.4]
  wire [15:0] _T_96843; // @[Mux.scala 31:69:@41249.4]
  wire [15:0] _T_96844; // @[Mux.scala 31:69:@41250.4]
  wire [15:0] _T_96845; // @[Mux.scala 31:69:@41251.4]
  wire  _T_96846; // @[OneHot.scala 66:30:@41252.4]
  wire  _T_96847; // @[OneHot.scala 66:30:@41253.4]
  wire  _T_96848; // @[OneHot.scala 66:30:@41254.4]
  wire  _T_96849; // @[OneHot.scala 66:30:@41255.4]
  wire  _T_96850; // @[OneHot.scala 66:30:@41256.4]
  wire  _T_96851; // @[OneHot.scala 66:30:@41257.4]
  wire  _T_96852; // @[OneHot.scala 66:30:@41258.4]
  wire  _T_96853; // @[OneHot.scala 66:30:@41259.4]
  wire  _T_96854; // @[OneHot.scala 66:30:@41260.4]
  wire  _T_96855; // @[OneHot.scala 66:30:@41261.4]
  wire  _T_96856; // @[OneHot.scala 66:30:@41262.4]
  wire  _T_96857; // @[OneHot.scala 66:30:@41263.4]
  wire  _T_96858; // @[OneHot.scala 66:30:@41264.4]
  wire  _T_96859; // @[OneHot.scala 66:30:@41265.4]
  wire  _T_96860; // @[OneHot.scala 66:30:@41266.4]
  wire  _T_96861; // @[OneHot.scala 66:30:@41267.4]
  wire [15:0] _T_96902; // @[Mux.scala 31:69:@41285.4]
  wire [15:0] _T_96903; // @[Mux.scala 31:69:@41286.4]
  wire [15:0] _T_96904; // @[Mux.scala 31:69:@41287.4]
  wire [15:0] _T_96905; // @[Mux.scala 31:69:@41288.4]
  wire [15:0] _T_96906; // @[Mux.scala 31:69:@41289.4]
  wire [15:0] _T_96907; // @[Mux.scala 31:69:@41290.4]
  wire [15:0] _T_96908; // @[Mux.scala 31:69:@41291.4]
  wire [15:0] _T_96909; // @[Mux.scala 31:69:@41292.4]
  wire [15:0] _T_96910; // @[Mux.scala 31:69:@41293.4]
  wire [15:0] _T_96911; // @[Mux.scala 31:69:@41294.4]
  wire [15:0] _T_96912; // @[Mux.scala 31:69:@41295.4]
  wire [15:0] _T_96913; // @[Mux.scala 31:69:@41296.4]
  wire [15:0] _T_96914; // @[Mux.scala 31:69:@41297.4]
  wire [15:0] _T_96915; // @[Mux.scala 31:69:@41298.4]
  wire [15:0] _T_96916; // @[Mux.scala 31:69:@41299.4]
  wire [15:0] _T_96917; // @[Mux.scala 31:69:@41300.4]
  wire  _T_96918; // @[OneHot.scala 66:30:@41301.4]
  wire  _T_96919; // @[OneHot.scala 66:30:@41302.4]
  wire  _T_96920; // @[OneHot.scala 66:30:@41303.4]
  wire  _T_96921; // @[OneHot.scala 66:30:@41304.4]
  wire  _T_96922; // @[OneHot.scala 66:30:@41305.4]
  wire  _T_96923; // @[OneHot.scala 66:30:@41306.4]
  wire  _T_96924; // @[OneHot.scala 66:30:@41307.4]
  wire  _T_96925; // @[OneHot.scala 66:30:@41308.4]
  wire  _T_96926; // @[OneHot.scala 66:30:@41309.4]
  wire  _T_96927; // @[OneHot.scala 66:30:@41310.4]
  wire  _T_96928; // @[OneHot.scala 66:30:@41311.4]
  wire  _T_96929; // @[OneHot.scala 66:30:@41312.4]
  wire  _T_96930; // @[OneHot.scala 66:30:@41313.4]
  wire  _T_96931; // @[OneHot.scala 66:30:@41314.4]
  wire  _T_96932; // @[OneHot.scala 66:30:@41315.4]
  wire  _T_96933; // @[OneHot.scala 66:30:@41316.4]
  wire [15:0] _T_96974; // @[Mux.scala 31:69:@41334.4]
  wire [15:0] _T_96975; // @[Mux.scala 31:69:@41335.4]
  wire [15:0] _T_96976; // @[Mux.scala 31:69:@41336.4]
  wire [15:0] _T_96977; // @[Mux.scala 31:69:@41337.4]
  wire [15:0] _T_96978; // @[Mux.scala 31:69:@41338.4]
  wire [15:0] _T_96979; // @[Mux.scala 31:69:@41339.4]
  wire [15:0] _T_96980; // @[Mux.scala 31:69:@41340.4]
  wire [15:0] _T_96981; // @[Mux.scala 31:69:@41341.4]
  wire [15:0] _T_96982; // @[Mux.scala 31:69:@41342.4]
  wire [15:0] _T_96983; // @[Mux.scala 31:69:@41343.4]
  wire [15:0] _T_96984; // @[Mux.scala 31:69:@41344.4]
  wire [15:0] _T_96985; // @[Mux.scala 31:69:@41345.4]
  wire [15:0] _T_96986; // @[Mux.scala 31:69:@41346.4]
  wire [15:0] _T_96987; // @[Mux.scala 31:69:@41347.4]
  wire [15:0] _T_96988; // @[Mux.scala 31:69:@41348.4]
  wire [15:0] _T_96989; // @[Mux.scala 31:69:@41349.4]
  wire  _T_96990; // @[OneHot.scala 66:30:@41350.4]
  wire  _T_96991; // @[OneHot.scala 66:30:@41351.4]
  wire  _T_96992; // @[OneHot.scala 66:30:@41352.4]
  wire  _T_96993; // @[OneHot.scala 66:30:@41353.4]
  wire  _T_96994; // @[OneHot.scala 66:30:@41354.4]
  wire  _T_96995; // @[OneHot.scala 66:30:@41355.4]
  wire  _T_96996; // @[OneHot.scala 66:30:@41356.4]
  wire  _T_96997; // @[OneHot.scala 66:30:@41357.4]
  wire  _T_96998; // @[OneHot.scala 66:30:@41358.4]
  wire  _T_96999; // @[OneHot.scala 66:30:@41359.4]
  wire  _T_97000; // @[OneHot.scala 66:30:@41360.4]
  wire  _T_97001; // @[OneHot.scala 66:30:@41361.4]
  wire  _T_97002; // @[OneHot.scala 66:30:@41362.4]
  wire  _T_97003; // @[OneHot.scala 66:30:@41363.4]
  wire  _T_97004; // @[OneHot.scala 66:30:@41364.4]
  wire  _T_97005; // @[OneHot.scala 66:30:@41365.4]
  wire [15:0] _T_97046; // @[Mux.scala 31:69:@41383.4]
  wire [15:0] _T_97047; // @[Mux.scala 31:69:@41384.4]
  wire [15:0] _T_97048; // @[Mux.scala 31:69:@41385.4]
  wire [15:0] _T_97049; // @[Mux.scala 31:69:@41386.4]
  wire [15:0] _T_97050; // @[Mux.scala 31:69:@41387.4]
  wire [15:0] _T_97051; // @[Mux.scala 31:69:@41388.4]
  wire [15:0] _T_97052; // @[Mux.scala 31:69:@41389.4]
  wire [15:0] _T_97053; // @[Mux.scala 31:69:@41390.4]
  wire [15:0] _T_97054; // @[Mux.scala 31:69:@41391.4]
  wire [15:0] _T_97055; // @[Mux.scala 31:69:@41392.4]
  wire [15:0] _T_97056; // @[Mux.scala 31:69:@41393.4]
  wire [15:0] _T_97057; // @[Mux.scala 31:69:@41394.4]
  wire [15:0] _T_97058; // @[Mux.scala 31:69:@41395.4]
  wire [15:0] _T_97059; // @[Mux.scala 31:69:@41396.4]
  wire [15:0] _T_97060; // @[Mux.scala 31:69:@41397.4]
  wire [15:0] _T_97061; // @[Mux.scala 31:69:@41398.4]
  wire  _T_97062; // @[OneHot.scala 66:30:@41399.4]
  wire  _T_97063; // @[OneHot.scala 66:30:@41400.4]
  wire  _T_97064; // @[OneHot.scala 66:30:@41401.4]
  wire  _T_97065; // @[OneHot.scala 66:30:@41402.4]
  wire  _T_97066; // @[OneHot.scala 66:30:@41403.4]
  wire  _T_97067; // @[OneHot.scala 66:30:@41404.4]
  wire  _T_97068; // @[OneHot.scala 66:30:@41405.4]
  wire  _T_97069; // @[OneHot.scala 66:30:@41406.4]
  wire  _T_97070; // @[OneHot.scala 66:30:@41407.4]
  wire  _T_97071; // @[OneHot.scala 66:30:@41408.4]
  wire  _T_97072; // @[OneHot.scala 66:30:@41409.4]
  wire  _T_97073; // @[OneHot.scala 66:30:@41410.4]
  wire  _T_97074; // @[OneHot.scala 66:30:@41411.4]
  wire  _T_97075; // @[OneHot.scala 66:30:@41412.4]
  wire  _T_97076; // @[OneHot.scala 66:30:@41413.4]
  wire  _T_97077; // @[OneHot.scala 66:30:@41414.4]
  wire [7:0] _T_97142; // @[Mux.scala 19:72:@41438.4]
  wire [15:0] _T_97150; // @[Mux.scala 19:72:@41446.4]
  wire [15:0] _T_97152; // @[Mux.scala 19:72:@41447.4]
  wire [7:0] _T_97159; // @[Mux.scala 19:72:@41454.4]
  wire [15:0] _T_97167; // @[Mux.scala 19:72:@41462.4]
  wire [15:0] _T_97169; // @[Mux.scala 19:72:@41463.4]
  wire [7:0] _T_97176; // @[Mux.scala 19:72:@41470.4]
  wire [15:0] _T_97184; // @[Mux.scala 19:72:@41478.4]
  wire [15:0] _T_97186; // @[Mux.scala 19:72:@41479.4]
  wire [7:0] _T_97193; // @[Mux.scala 19:72:@41486.4]
  wire [15:0] _T_97201; // @[Mux.scala 19:72:@41494.4]
  wire [15:0] _T_97203; // @[Mux.scala 19:72:@41495.4]
  wire [7:0] _T_97210; // @[Mux.scala 19:72:@41502.4]
  wire [15:0] _T_97218; // @[Mux.scala 19:72:@41510.4]
  wire [15:0] _T_97220; // @[Mux.scala 19:72:@41511.4]
  wire [7:0] _T_97227; // @[Mux.scala 19:72:@41518.4]
  wire [15:0] _T_97235; // @[Mux.scala 19:72:@41526.4]
  wire [15:0] _T_97237; // @[Mux.scala 19:72:@41527.4]
  wire [7:0] _T_97244; // @[Mux.scala 19:72:@41534.4]
  wire [15:0] _T_97252; // @[Mux.scala 19:72:@41542.4]
  wire [15:0] _T_97254; // @[Mux.scala 19:72:@41543.4]
  wire [7:0] _T_97261; // @[Mux.scala 19:72:@41550.4]
  wire [15:0] _T_97269; // @[Mux.scala 19:72:@41558.4]
  wire [15:0] _T_97271; // @[Mux.scala 19:72:@41559.4]
  wire [7:0] _T_97278; // @[Mux.scala 19:72:@41566.4]
  wire [15:0] _T_97286; // @[Mux.scala 19:72:@41574.4]
  wire [15:0] _T_97288; // @[Mux.scala 19:72:@41575.4]
  wire [7:0] _T_97295; // @[Mux.scala 19:72:@41582.4]
  wire [15:0] _T_97303; // @[Mux.scala 19:72:@41590.4]
  wire [15:0] _T_97305; // @[Mux.scala 19:72:@41591.4]
  wire [7:0] _T_97312; // @[Mux.scala 19:72:@41598.4]
  wire [15:0] _T_97320; // @[Mux.scala 19:72:@41606.4]
  wire [15:0] _T_97322; // @[Mux.scala 19:72:@41607.4]
  wire [7:0] _T_97329; // @[Mux.scala 19:72:@41614.4]
  wire [15:0] _T_97337; // @[Mux.scala 19:72:@41622.4]
  wire [15:0] _T_97339; // @[Mux.scala 19:72:@41623.4]
  wire [7:0] _T_97346; // @[Mux.scala 19:72:@41630.4]
  wire [15:0] _T_97354; // @[Mux.scala 19:72:@41638.4]
  wire [15:0] _T_97356; // @[Mux.scala 19:72:@41639.4]
  wire [7:0] _T_97363; // @[Mux.scala 19:72:@41646.4]
  wire [15:0] _T_97371; // @[Mux.scala 19:72:@41654.4]
  wire [15:0] _T_97373; // @[Mux.scala 19:72:@41655.4]
  wire [7:0] _T_97380; // @[Mux.scala 19:72:@41662.4]
  wire [15:0] _T_97388; // @[Mux.scala 19:72:@41670.4]
  wire [15:0] _T_97390; // @[Mux.scala 19:72:@41671.4]
  wire [7:0] _T_97397; // @[Mux.scala 19:72:@41678.4]
  wire [15:0] _T_97405; // @[Mux.scala 19:72:@41686.4]
  wire [15:0] _T_97407; // @[Mux.scala 19:72:@41687.4]
  wire [15:0] _T_97408; // @[Mux.scala 19:72:@41688.4]
  wire [15:0] _T_97409; // @[Mux.scala 19:72:@41689.4]
  wire [15:0] _T_97410; // @[Mux.scala 19:72:@41690.4]
  wire [15:0] _T_97411; // @[Mux.scala 19:72:@41691.4]
  wire [15:0] _T_97412; // @[Mux.scala 19:72:@41692.4]
  wire [15:0] _T_97413; // @[Mux.scala 19:72:@41693.4]
  wire [15:0] _T_97414; // @[Mux.scala 19:72:@41694.4]
  wire [15:0] _T_97415; // @[Mux.scala 19:72:@41695.4]
  wire [15:0] _T_97416; // @[Mux.scala 19:72:@41696.4]
  wire [15:0] _T_97417; // @[Mux.scala 19:72:@41697.4]
  wire [15:0] _T_97418; // @[Mux.scala 19:72:@41698.4]
  wire [15:0] _T_97419; // @[Mux.scala 19:72:@41699.4]
  wire [15:0] _T_97420; // @[Mux.scala 19:72:@41700.4]
  wire [15:0] _T_97421; // @[Mux.scala 19:72:@41701.4]
  wire [15:0] _T_97422; // @[Mux.scala 19:72:@41702.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@41706.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@41708.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@41710.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@41712.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@41714.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@41716.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@41718.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@41720.4]
  wire  outputPriorityPorts_0_8; // @[Mux.scala 19:72:@41722.4]
  wire  outputPriorityPorts_0_9; // @[Mux.scala 19:72:@41724.4]
  wire  outputPriorityPorts_0_10; // @[Mux.scala 19:72:@41726.4]
  wire  outputPriorityPorts_0_11; // @[Mux.scala 19:72:@41728.4]
  wire  outputPriorityPorts_0_12; // @[Mux.scala 19:72:@41730.4]
  wire  outputPriorityPorts_0_13; // @[Mux.scala 19:72:@41732.4]
  wire  outputPriorityPorts_0_14; // @[Mux.scala 19:72:@41734.4]
  wire  outputPriorityPorts_0_15; // @[Mux.scala 19:72:@41736.4]
  wire  _T_97565; // @[LoadQueue.scala 313:47:@41758.6]
  wire [31:0] _GEN_2114; // @[LoadQueue.scala 314:36:@41762.6]
  wire  _GEN_2115; // @[LoadQueue.scala 314:36:@41762.6]
  wire  _GEN_2116; // @[LoadQueue.scala 308:34:@41754.4]
  wire [31:0] _GEN_2117; // @[LoadQueue.scala 308:34:@41754.4]
  wire  _T_97580; // @[LoadQueue.scala 313:47:@41771.6]
  wire [31:0] _GEN_2118; // @[LoadQueue.scala 314:36:@41775.6]
  wire  _GEN_2119; // @[LoadQueue.scala 314:36:@41775.6]
  wire  _GEN_2120; // @[LoadQueue.scala 308:34:@41767.4]
  wire [31:0] _GEN_2121; // @[LoadQueue.scala 308:34:@41767.4]
  wire  _T_97595; // @[LoadQueue.scala 313:47:@41784.6]
  wire [31:0] _GEN_2122; // @[LoadQueue.scala 314:36:@41788.6]
  wire  _GEN_2123; // @[LoadQueue.scala 314:36:@41788.6]
  wire  _GEN_2124; // @[LoadQueue.scala 308:34:@41780.4]
  wire [31:0] _GEN_2125; // @[LoadQueue.scala 308:34:@41780.4]
  wire  _T_97610; // @[LoadQueue.scala 313:47:@41797.6]
  wire [31:0] _GEN_2126; // @[LoadQueue.scala 314:36:@41801.6]
  wire  _GEN_2127; // @[LoadQueue.scala 314:36:@41801.6]
  wire  _GEN_2128; // @[LoadQueue.scala 308:34:@41793.4]
  wire [31:0] _GEN_2129; // @[LoadQueue.scala 308:34:@41793.4]
  wire  _T_97625; // @[LoadQueue.scala 313:47:@41810.6]
  wire [31:0] _GEN_2130; // @[LoadQueue.scala 314:36:@41814.6]
  wire  _GEN_2131; // @[LoadQueue.scala 314:36:@41814.6]
  wire  _GEN_2132; // @[LoadQueue.scala 308:34:@41806.4]
  wire [31:0] _GEN_2133; // @[LoadQueue.scala 308:34:@41806.4]
  wire  _T_97640; // @[LoadQueue.scala 313:47:@41823.6]
  wire [31:0] _GEN_2134; // @[LoadQueue.scala 314:36:@41827.6]
  wire  _GEN_2135; // @[LoadQueue.scala 314:36:@41827.6]
  wire  _GEN_2136; // @[LoadQueue.scala 308:34:@41819.4]
  wire [31:0] _GEN_2137; // @[LoadQueue.scala 308:34:@41819.4]
  wire  _T_97655; // @[LoadQueue.scala 313:47:@41836.6]
  wire [31:0] _GEN_2138; // @[LoadQueue.scala 314:36:@41840.6]
  wire  _GEN_2139; // @[LoadQueue.scala 314:36:@41840.6]
  wire  _GEN_2140; // @[LoadQueue.scala 308:34:@41832.4]
  wire [31:0] _GEN_2141; // @[LoadQueue.scala 308:34:@41832.4]
  wire  _T_97670; // @[LoadQueue.scala 313:47:@41849.6]
  wire [31:0] _GEN_2142; // @[LoadQueue.scala 314:36:@41853.6]
  wire  _GEN_2143; // @[LoadQueue.scala 314:36:@41853.6]
  wire  _GEN_2144; // @[LoadQueue.scala 308:34:@41845.4]
  wire [31:0] _GEN_2145; // @[LoadQueue.scala 308:34:@41845.4]
  wire  _T_97685; // @[LoadQueue.scala 313:47:@41862.6]
  wire [31:0] _GEN_2146; // @[LoadQueue.scala 314:36:@41866.6]
  wire  _GEN_2147; // @[LoadQueue.scala 314:36:@41866.6]
  wire  _GEN_2148; // @[LoadQueue.scala 308:34:@41858.4]
  wire [31:0] _GEN_2149; // @[LoadQueue.scala 308:34:@41858.4]
  wire  _T_97700; // @[LoadQueue.scala 313:47:@41875.6]
  wire [31:0] _GEN_2150; // @[LoadQueue.scala 314:36:@41879.6]
  wire  _GEN_2151; // @[LoadQueue.scala 314:36:@41879.6]
  wire  _GEN_2152; // @[LoadQueue.scala 308:34:@41871.4]
  wire [31:0] _GEN_2153; // @[LoadQueue.scala 308:34:@41871.4]
  wire  _T_97715; // @[LoadQueue.scala 313:47:@41888.6]
  wire [31:0] _GEN_2154; // @[LoadQueue.scala 314:36:@41892.6]
  wire  _GEN_2155; // @[LoadQueue.scala 314:36:@41892.6]
  wire  _GEN_2156; // @[LoadQueue.scala 308:34:@41884.4]
  wire [31:0] _GEN_2157; // @[LoadQueue.scala 308:34:@41884.4]
  wire  _T_97730; // @[LoadQueue.scala 313:47:@41901.6]
  wire [31:0] _GEN_2158; // @[LoadQueue.scala 314:36:@41905.6]
  wire  _GEN_2159; // @[LoadQueue.scala 314:36:@41905.6]
  wire  _GEN_2160; // @[LoadQueue.scala 308:34:@41897.4]
  wire [31:0] _GEN_2161; // @[LoadQueue.scala 308:34:@41897.4]
  wire  _T_97745; // @[LoadQueue.scala 313:47:@41914.6]
  wire [31:0] _GEN_2162; // @[LoadQueue.scala 314:36:@41918.6]
  wire  _GEN_2163; // @[LoadQueue.scala 314:36:@41918.6]
  wire  _GEN_2164; // @[LoadQueue.scala 308:34:@41910.4]
  wire [31:0] _GEN_2165; // @[LoadQueue.scala 308:34:@41910.4]
  wire  _T_97760; // @[LoadQueue.scala 313:47:@41927.6]
  wire [31:0] _GEN_2166; // @[LoadQueue.scala 314:36:@41931.6]
  wire  _GEN_2167; // @[LoadQueue.scala 314:36:@41931.6]
  wire  _GEN_2168; // @[LoadQueue.scala 308:34:@41923.4]
  wire [31:0] _GEN_2169; // @[LoadQueue.scala 308:34:@41923.4]
  wire  _T_97775; // @[LoadQueue.scala 313:47:@41940.6]
  wire [31:0] _GEN_2170; // @[LoadQueue.scala 314:36:@41944.6]
  wire  _GEN_2171; // @[LoadQueue.scala 314:36:@41944.6]
  wire  _GEN_2172; // @[LoadQueue.scala 308:34:@41936.4]
  wire [31:0] _GEN_2173; // @[LoadQueue.scala 308:34:@41936.4]
  wire  _T_97790; // @[LoadQueue.scala 313:47:@41953.6]
  wire [31:0] _GEN_2174; // @[LoadQueue.scala 314:36:@41957.6]
  wire  _GEN_2175; // @[LoadQueue.scala 314:36:@41957.6]
  wire  _GEN_2176; // @[LoadQueue.scala 308:34:@41949.4]
  wire [31:0] _GEN_2177; // @[LoadQueue.scala 308:34:@41949.4]
  wire  _T_97825; // @[LoadQueue.scala 326:108:@41963.4]
  wire  _T_97827; // @[LoadQueue.scala 327:34:@41964.4]
  wire  _T_97828; // @[LoadQueue.scala 327:31:@41965.4]
  wire  loadCompleting_0; // @[LoadQueue.scala 327:63:@41966.4]
  wire  _T_97839; // @[LoadQueue.scala 326:108:@41971.4]
  wire  _T_97841; // @[LoadQueue.scala 327:34:@41972.4]
  wire  _T_97842; // @[LoadQueue.scala 327:31:@41973.4]
  wire  loadCompleting_1; // @[LoadQueue.scala 327:63:@41974.4]
  wire  _T_97853; // @[LoadQueue.scala 326:108:@41979.4]
  wire  _T_97855; // @[LoadQueue.scala 327:34:@41980.4]
  wire  _T_97856; // @[LoadQueue.scala 327:31:@41981.4]
  wire  loadCompleting_2; // @[LoadQueue.scala 327:63:@41982.4]
  wire  _T_97867; // @[LoadQueue.scala 326:108:@41987.4]
  wire  _T_97869; // @[LoadQueue.scala 327:34:@41988.4]
  wire  _T_97870; // @[LoadQueue.scala 327:31:@41989.4]
  wire  loadCompleting_3; // @[LoadQueue.scala 327:63:@41990.4]
  wire  _T_97881; // @[LoadQueue.scala 326:108:@41995.4]
  wire  _T_97883; // @[LoadQueue.scala 327:34:@41996.4]
  wire  _T_97884; // @[LoadQueue.scala 327:31:@41997.4]
  wire  loadCompleting_4; // @[LoadQueue.scala 327:63:@41998.4]
  wire  _T_97895; // @[LoadQueue.scala 326:108:@42003.4]
  wire  _T_97897; // @[LoadQueue.scala 327:34:@42004.4]
  wire  _T_97898; // @[LoadQueue.scala 327:31:@42005.4]
  wire  loadCompleting_5; // @[LoadQueue.scala 327:63:@42006.4]
  wire  _T_97909; // @[LoadQueue.scala 326:108:@42011.4]
  wire  _T_97911; // @[LoadQueue.scala 327:34:@42012.4]
  wire  _T_97912; // @[LoadQueue.scala 327:31:@42013.4]
  wire  loadCompleting_6; // @[LoadQueue.scala 327:63:@42014.4]
  wire  _T_97923; // @[LoadQueue.scala 326:108:@42019.4]
  wire  _T_97925; // @[LoadQueue.scala 327:34:@42020.4]
  wire  _T_97926; // @[LoadQueue.scala 327:31:@42021.4]
  wire  loadCompleting_7; // @[LoadQueue.scala 327:63:@42022.4]
  wire  _T_97937; // @[LoadQueue.scala 326:108:@42027.4]
  wire  _T_97939; // @[LoadQueue.scala 327:34:@42028.4]
  wire  _T_97940; // @[LoadQueue.scala 327:31:@42029.4]
  wire  loadCompleting_8; // @[LoadQueue.scala 327:63:@42030.4]
  wire  _T_97951; // @[LoadQueue.scala 326:108:@42035.4]
  wire  _T_97953; // @[LoadQueue.scala 327:34:@42036.4]
  wire  _T_97954; // @[LoadQueue.scala 327:31:@42037.4]
  wire  loadCompleting_9; // @[LoadQueue.scala 327:63:@42038.4]
  wire  _T_97965; // @[LoadQueue.scala 326:108:@42043.4]
  wire  _T_97967; // @[LoadQueue.scala 327:34:@42044.4]
  wire  _T_97968; // @[LoadQueue.scala 327:31:@42045.4]
  wire  loadCompleting_10; // @[LoadQueue.scala 327:63:@42046.4]
  wire  _T_97979; // @[LoadQueue.scala 326:108:@42051.4]
  wire  _T_97981; // @[LoadQueue.scala 327:34:@42052.4]
  wire  _T_97982; // @[LoadQueue.scala 327:31:@42053.4]
  wire  loadCompleting_11; // @[LoadQueue.scala 327:63:@42054.4]
  wire  _T_97993; // @[LoadQueue.scala 326:108:@42059.4]
  wire  _T_97995; // @[LoadQueue.scala 327:34:@42060.4]
  wire  _T_97996; // @[LoadQueue.scala 327:31:@42061.4]
  wire  loadCompleting_12; // @[LoadQueue.scala 327:63:@42062.4]
  wire  _T_98007; // @[LoadQueue.scala 326:108:@42067.4]
  wire  _T_98009; // @[LoadQueue.scala 327:34:@42068.4]
  wire  _T_98010; // @[LoadQueue.scala 327:31:@42069.4]
  wire  loadCompleting_13; // @[LoadQueue.scala 327:63:@42070.4]
  wire  _T_98021; // @[LoadQueue.scala 326:108:@42075.4]
  wire  _T_98023; // @[LoadQueue.scala 327:34:@42076.4]
  wire  _T_98024; // @[LoadQueue.scala 327:31:@42077.4]
  wire  loadCompleting_14; // @[LoadQueue.scala 327:63:@42078.4]
  wire  _T_98035; // @[LoadQueue.scala 326:108:@42083.4]
  wire  _T_98037; // @[LoadQueue.scala 327:34:@42084.4]
  wire  _T_98038; // @[LoadQueue.scala 327:31:@42085.4]
  wire  loadCompleting_15; // @[LoadQueue.scala 327:63:@42086.4]
  wire  _GEN_2178; // @[LoadQueue.scala 337:46:@42095.6]
  wire  _GEN_2179; // @[LoadQueue.scala 335:34:@42091.4]
  wire  _GEN_2180; // @[LoadQueue.scala 337:46:@42102.6]
  wire  _GEN_2181; // @[LoadQueue.scala 335:34:@42098.4]
  wire  _GEN_2182; // @[LoadQueue.scala 337:46:@42109.6]
  wire  _GEN_2183; // @[LoadQueue.scala 335:34:@42105.4]
  wire  _GEN_2184; // @[LoadQueue.scala 337:46:@42116.6]
  wire  _GEN_2185; // @[LoadQueue.scala 335:34:@42112.4]
  wire  _GEN_2186; // @[LoadQueue.scala 337:46:@42123.6]
  wire  _GEN_2187; // @[LoadQueue.scala 335:34:@42119.4]
  wire  _GEN_2188; // @[LoadQueue.scala 337:46:@42130.6]
  wire  _GEN_2189; // @[LoadQueue.scala 335:34:@42126.4]
  wire  _GEN_2190; // @[LoadQueue.scala 337:46:@42137.6]
  wire  _GEN_2191; // @[LoadQueue.scala 335:34:@42133.4]
  wire  _GEN_2192; // @[LoadQueue.scala 337:46:@42144.6]
  wire  _GEN_2193; // @[LoadQueue.scala 335:34:@42140.4]
  wire  _GEN_2194; // @[LoadQueue.scala 337:46:@42151.6]
  wire  _GEN_2195; // @[LoadQueue.scala 335:34:@42147.4]
  wire  _GEN_2196; // @[LoadQueue.scala 337:46:@42158.6]
  wire  _GEN_2197; // @[LoadQueue.scala 335:34:@42154.4]
  wire  _GEN_2198; // @[LoadQueue.scala 337:46:@42165.6]
  wire  _GEN_2199; // @[LoadQueue.scala 335:34:@42161.4]
  wire  _GEN_2200; // @[LoadQueue.scala 337:46:@42172.6]
  wire  _GEN_2201; // @[LoadQueue.scala 335:34:@42168.4]
  wire  _GEN_2202; // @[LoadQueue.scala 337:46:@42179.6]
  wire  _GEN_2203; // @[LoadQueue.scala 335:34:@42175.4]
  wire  _GEN_2204; // @[LoadQueue.scala 337:46:@42186.6]
  wire  _GEN_2205; // @[LoadQueue.scala 335:34:@42182.4]
  wire  _GEN_2206; // @[LoadQueue.scala 337:46:@42193.6]
  wire  _GEN_2207; // @[LoadQueue.scala 335:34:@42189.4]
  wire  _GEN_2208; // @[LoadQueue.scala 337:46:@42200.6]
  wire  _GEN_2209; // @[LoadQueue.scala 335:34:@42196.4]
  wire  _T_98169; // @[LoadQueue.scala 348:24:@42269.4]
  wire  _T_98170; // @[LoadQueue.scala 348:24:@42270.4]
  wire  _T_98171; // @[LoadQueue.scala 348:24:@42271.4]
  wire  _T_98172; // @[LoadQueue.scala 348:24:@42272.4]
  wire  _T_98173; // @[LoadQueue.scala 348:24:@42273.4]
  wire  _T_98174; // @[LoadQueue.scala 348:24:@42274.4]
  wire  _T_98175; // @[LoadQueue.scala 348:24:@42275.4]
  wire  _T_98176; // @[LoadQueue.scala 348:24:@42276.4]
  wire  _T_98177; // @[LoadQueue.scala 348:24:@42277.4]
  wire  _T_98178; // @[LoadQueue.scala 348:24:@42278.4]
  wire  _T_98179; // @[LoadQueue.scala 348:24:@42279.4]
  wire  _T_98180; // @[LoadQueue.scala 348:24:@42280.4]
  wire  _T_98181; // @[LoadQueue.scala 348:24:@42281.4]
  wire  _T_98182; // @[LoadQueue.scala 348:24:@42282.4]
  wire  _T_98183; // @[LoadQueue.scala 348:24:@42283.4]
  wire [3:0] _T_98200; // @[Mux.scala 31:69:@42285.6]
  wire [3:0] _T_98201; // @[Mux.scala 31:69:@42286.6]
  wire [3:0] _T_98202; // @[Mux.scala 31:69:@42287.6]
  wire [3:0] _T_98203; // @[Mux.scala 31:69:@42288.6]
  wire [3:0] _T_98204; // @[Mux.scala 31:69:@42289.6]
  wire [3:0] _T_98205; // @[Mux.scala 31:69:@42290.6]
  wire [3:0] _T_98206; // @[Mux.scala 31:69:@42291.6]
  wire [3:0] _T_98207; // @[Mux.scala 31:69:@42292.6]
  wire [3:0] _T_98208; // @[Mux.scala 31:69:@42293.6]
  wire [3:0] _T_98209; // @[Mux.scala 31:69:@42294.6]
  wire [3:0] _T_98210; // @[Mux.scala 31:69:@42295.6]
  wire [3:0] _T_98211; // @[Mux.scala 31:69:@42296.6]
  wire [3:0] _T_98212; // @[Mux.scala 31:69:@42297.6]
  wire [3:0] _T_98213; // @[Mux.scala 31:69:@42298.6]
  wire [3:0] _T_98214; // @[Mux.scala 31:69:@42299.6]
  wire [31:0] _GEN_2211; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2212; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2213; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2214; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2215; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2216; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2217; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2218; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2219; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2220; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2221; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2222; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2223; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2224; // @[LoadQueue.scala 349:37:@42300.6]
  wire [31:0] _GEN_2225; // @[LoadQueue.scala 349:37:@42300.6]
  wire  _GEN_2229; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2230; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2231; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2232; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2233; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2234; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2235; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2236; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2237; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2238; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2239; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2240; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2241; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2242; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2243; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2245; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2246; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2247; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2248; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2249; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2250; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2251; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2252; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2253; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2254; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2255; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2256; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2257; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2258; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _GEN_2259; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _T_98225; // @[LoadQueue.scala 363:29:@42307.4]
  wire  _T_98226; // @[LoadQueue.scala 363:63:@42308.4]
  wire  _T_98228; // @[LoadQueue.scala 363:75:@42309.4]
  wire  _T_98229; // @[LoadQueue.scala 363:72:@42310.4]
  wire  _T_98230; // @[LoadQueue.scala 363:54:@42311.4]
  wire [4:0] _T_98233; // @[util.scala 10:8:@42313.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@42314.6]
  wire [4:0] _T_98234; // @[util.scala 10:14:@42314.6]
  wire [4:0] _GEN_2260; // @[LoadQueue.scala 363:91:@42312.4]
  wire [3:0] _GEN_2358; // @[util.scala 10:8:@42318.6]
  wire [4:0] _T_98236; // @[util.scala 10:8:@42318.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@42319.6]
  wire [4:0] _T_98237; // @[util.scala 10:14:@42319.6]
  wire [4:0] _GEN_2261; // @[LoadQueue.scala 367:20:@42317.4]
  wire  _T_98239; // @[LoadQueue.scala 371:82:@42322.4]
  wire  _T_98240; // @[LoadQueue.scala 371:79:@42323.4]
  wire  _T_98242; // @[LoadQueue.scala 371:82:@42324.4]
  wire  _T_98243; // @[LoadQueue.scala 371:79:@42325.4]
  wire  _T_98245; // @[LoadQueue.scala 371:82:@42326.4]
  wire  _T_98246; // @[LoadQueue.scala 371:79:@42327.4]
  wire  _T_98248; // @[LoadQueue.scala 371:82:@42328.4]
  wire  _T_98249; // @[LoadQueue.scala 371:79:@42329.4]
  wire  _T_98251; // @[LoadQueue.scala 371:82:@42330.4]
  wire  _T_98252; // @[LoadQueue.scala 371:79:@42331.4]
  wire  _T_98254; // @[LoadQueue.scala 371:82:@42332.4]
  wire  _T_98255; // @[LoadQueue.scala 371:79:@42333.4]
  wire  _T_98257; // @[LoadQueue.scala 371:82:@42334.4]
  wire  _T_98258; // @[LoadQueue.scala 371:79:@42335.4]
  wire  _T_98260; // @[LoadQueue.scala 371:82:@42336.4]
  wire  _T_98261; // @[LoadQueue.scala 371:79:@42337.4]
  wire  _T_98263; // @[LoadQueue.scala 371:82:@42338.4]
  wire  _T_98264; // @[LoadQueue.scala 371:79:@42339.4]
  wire  _T_98266; // @[LoadQueue.scala 371:82:@42340.4]
  wire  _T_98267; // @[LoadQueue.scala 371:79:@42341.4]
  wire  _T_98269; // @[LoadQueue.scala 371:82:@42342.4]
  wire  _T_98270; // @[LoadQueue.scala 371:79:@42343.4]
  wire  _T_98272; // @[LoadQueue.scala 371:82:@42344.4]
  wire  _T_98273; // @[LoadQueue.scala 371:79:@42345.4]
  wire  _T_98275; // @[LoadQueue.scala 371:82:@42346.4]
  wire  _T_98276; // @[LoadQueue.scala 371:79:@42347.4]
  wire  _T_98278; // @[LoadQueue.scala 371:82:@42348.4]
  wire  _T_98279; // @[LoadQueue.scala 371:79:@42349.4]
  wire  _T_98281; // @[LoadQueue.scala 371:82:@42350.4]
  wire  _T_98282; // @[LoadQueue.scala 371:79:@42351.4]
  wire  _T_98284; // @[LoadQueue.scala 371:82:@42352.4]
  wire  _T_98285; // @[LoadQueue.scala 371:79:@42353.4]
  wire  _T_98310; // @[LoadQueue.scala 371:96:@42372.4]
  wire  _T_98311; // @[LoadQueue.scala 371:96:@42373.4]
  wire  _T_98312; // @[LoadQueue.scala 371:96:@42374.4]
  wire  _T_98313; // @[LoadQueue.scala 371:96:@42375.4]
  wire  _T_98314; // @[LoadQueue.scala 371:96:@42376.4]
  wire  _T_98315; // @[LoadQueue.scala 371:96:@42377.4]
  wire  _T_98316; // @[LoadQueue.scala 371:96:@42378.4]
  wire  _T_98317; // @[LoadQueue.scala 371:96:@42379.4]
  wire  _T_98318; // @[LoadQueue.scala 371:96:@42380.4]
  wire  _T_98319; // @[LoadQueue.scala 371:96:@42381.4]
  wire  _T_98320; // @[LoadQueue.scala 371:96:@42382.4]
  wire  _T_98321; // @[LoadQueue.scala 371:96:@42383.4]
  wire  _T_98322; // @[LoadQueue.scala 371:96:@42384.4]
  wire  _T_98323; // @[LoadQueue.scala 371:96:@42385.4]
  assign _GEN_2262 = {{2'd0}, tail}; // @[util.scala 14:20:@5032.4]
  assign _T_1716 = 6'h10 - _GEN_2262; // @[util.scala 14:20:@5032.4]
  assign _T_1717 = $unsigned(_T_1716); // @[util.scala 14:20:@5033.4]
  assign _T_1718 = _T_1717[5:0]; // @[util.scala 14:20:@5034.4]
  assign _GEN_0 = _T_1718 % 6'h10; // @[util.scala 14:25:@5035.4]
  assign _T_1719 = _GEN_0[4:0]; // @[util.scala 14:25:@5035.4]
  assign _GEN_2263 = {{4'd0}, io_bbNumLoads}; // @[LoadQueue.scala 71:46:@5036.4]
  assign _T_1720 = _T_1719 < _GEN_2263; // @[LoadQueue.scala 71:46:@5036.4]
  assign initBits_0 = _T_1720 & io_bbStart; // @[LoadQueue.scala 71:63:@5037.4]
  assign _T_1725 = 6'h11 - _GEN_2262; // @[util.scala 14:20:@5039.4]
  assign _T_1726 = $unsigned(_T_1725); // @[util.scala 14:20:@5040.4]
  assign _T_1727 = _T_1726[5:0]; // @[util.scala 14:20:@5041.4]
  assign _GEN_16 = _T_1727 % 6'h10; // @[util.scala 14:25:@5042.4]
  assign _T_1728 = _GEN_16[4:0]; // @[util.scala 14:25:@5042.4]
  assign _T_1729 = _T_1728 < _GEN_2263; // @[LoadQueue.scala 71:46:@5043.4]
  assign initBits_1 = _T_1729 & io_bbStart; // @[LoadQueue.scala 71:63:@5044.4]
  assign _T_1734 = 6'h12 - _GEN_2262; // @[util.scala 14:20:@5046.4]
  assign _T_1735 = $unsigned(_T_1734); // @[util.scala 14:20:@5047.4]
  assign _T_1736 = _T_1735[5:0]; // @[util.scala 14:20:@5048.4]
  assign _GEN_17 = _T_1736 % 6'h10; // @[util.scala 14:25:@5049.4]
  assign _T_1737 = _GEN_17[4:0]; // @[util.scala 14:25:@5049.4]
  assign _T_1738 = _T_1737 < _GEN_2263; // @[LoadQueue.scala 71:46:@5050.4]
  assign initBits_2 = _T_1738 & io_bbStart; // @[LoadQueue.scala 71:63:@5051.4]
  assign _T_1743 = 6'h13 - _GEN_2262; // @[util.scala 14:20:@5053.4]
  assign _T_1744 = $unsigned(_T_1743); // @[util.scala 14:20:@5054.4]
  assign _T_1745 = _T_1744[5:0]; // @[util.scala 14:20:@5055.4]
  assign _GEN_18 = _T_1745 % 6'h10; // @[util.scala 14:25:@5056.4]
  assign _T_1746 = _GEN_18[4:0]; // @[util.scala 14:25:@5056.4]
  assign _T_1747 = _T_1746 < _GEN_2263; // @[LoadQueue.scala 71:46:@5057.4]
  assign initBits_3 = _T_1747 & io_bbStart; // @[LoadQueue.scala 71:63:@5058.4]
  assign _T_1752 = 6'h14 - _GEN_2262; // @[util.scala 14:20:@5060.4]
  assign _T_1753 = $unsigned(_T_1752); // @[util.scala 14:20:@5061.4]
  assign _T_1754 = _T_1753[5:0]; // @[util.scala 14:20:@5062.4]
  assign _GEN_19 = _T_1754 % 6'h10; // @[util.scala 14:25:@5063.4]
  assign _T_1755 = _GEN_19[4:0]; // @[util.scala 14:25:@5063.4]
  assign _T_1756 = _T_1755 < _GEN_2263; // @[LoadQueue.scala 71:46:@5064.4]
  assign initBits_4 = _T_1756 & io_bbStart; // @[LoadQueue.scala 71:63:@5065.4]
  assign _T_1761 = 6'h15 - _GEN_2262; // @[util.scala 14:20:@5067.4]
  assign _T_1762 = $unsigned(_T_1761); // @[util.scala 14:20:@5068.4]
  assign _T_1763 = _T_1762[5:0]; // @[util.scala 14:20:@5069.4]
  assign _GEN_20 = _T_1763 % 6'h10; // @[util.scala 14:25:@5070.4]
  assign _T_1764 = _GEN_20[4:0]; // @[util.scala 14:25:@5070.4]
  assign _T_1765 = _T_1764 < _GEN_2263; // @[LoadQueue.scala 71:46:@5071.4]
  assign initBits_5 = _T_1765 & io_bbStart; // @[LoadQueue.scala 71:63:@5072.4]
  assign _T_1770 = 6'h16 - _GEN_2262; // @[util.scala 14:20:@5074.4]
  assign _T_1771 = $unsigned(_T_1770); // @[util.scala 14:20:@5075.4]
  assign _T_1772 = _T_1771[5:0]; // @[util.scala 14:20:@5076.4]
  assign _GEN_21 = _T_1772 % 6'h10; // @[util.scala 14:25:@5077.4]
  assign _T_1773 = _GEN_21[4:0]; // @[util.scala 14:25:@5077.4]
  assign _T_1774 = _T_1773 < _GEN_2263; // @[LoadQueue.scala 71:46:@5078.4]
  assign initBits_6 = _T_1774 & io_bbStart; // @[LoadQueue.scala 71:63:@5079.4]
  assign _T_1779 = 6'h17 - _GEN_2262; // @[util.scala 14:20:@5081.4]
  assign _T_1780 = $unsigned(_T_1779); // @[util.scala 14:20:@5082.4]
  assign _T_1781 = _T_1780[5:0]; // @[util.scala 14:20:@5083.4]
  assign _GEN_22 = _T_1781 % 6'h10; // @[util.scala 14:25:@5084.4]
  assign _T_1782 = _GEN_22[4:0]; // @[util.scala 14:25:@5084.4]
  assign _T_1783 = _T_1782 < _GEN_2263; // @[LoadQueue.scala 71:46:@5085.4]
  assign initBits_7 = _T_1783 & io_bbStart; // @[LoadQueue.scala 71:63:@5086.4]
  assign _T_1788 = 6'h18 - _GEN_2262; // @[util.scala 14:20:@5088.4]
  assign _T_1789 = $unsigned(_T_1788); // @[util.scala 14:20:@5089.4]
  assign _T_1790 = _T_1789[5:0]; // @[util.scala 14:20:@5090.4]
  assign _GEN_23 = _T_1790 % 6'h10; // @[util.scala 14:25:@5091.4]
  assign _T_1791 = _GEN_23[4:0]; // @[util.scala 14:25:@5091.4]
  assign _T_1792 = _T_1791 < _GEN_2263; // @[LoadQueue.scala 71:46:@5092.4]
  assign initBits_8 = _T_1792 & io_bbStart; // @[LoadQueue.scala 71:63:@5093.4]
  assign _T_1797 = 6'h19 - _GEN_2262; // @[util.scala 14:20:@5095.4]
  assign _T_1798 = $unsigned(_T_1797); // @[util.scala 14:20:@5096.4]
  assign _T_1799 = _T_1798[5:0]; // @[util.scala 14:20:@5097.4]
  assign _GEN_24 = _T_1799 % 6'h10; // @[util.scala 14:25:@5098.4]
  assign _T_1800 = _GEN_24[4:0]; // @[util.scala 14:25:@5098.4]
  assign _T_1801 = _T_1800 < _GEN_2263; // @[LoadQueue.scala 71:46:@5099.4]
  assign initBits_9 = _T_1801 & io_bbStart; // @[LoadQueue.scala 71:63:@5100.4]
  assign _T_1806 = 6'h1a - _GEN_2262; // @[util.scala 14:20:@5102.4]
  assign _T_1807 = $unsigned(_T_1806); // @[util.scala 14:20:@5103.4]
  assign _T_1808 = _T_1807[5:0]; // @[util.scala 14:20:@5104.4]
  assign _GEN_25 = _T_1808 % 6'h10; // @[util.scala 14:25:@5105.4]
  assign _T_1809 = _GEN_25[4:0]; // @[util.scala 14:25:@5105.4]
  assign _T_1810 = _T_1809 < _GEN_2263; // @[LoadQueue.scala 71:46:@5106.4]
  assign initBits_10 = _T_1810 & io_bbStart; // @[LoadQueue.scala 71:63:@5107.4]
  assign _T_1815 = 6'h1b - _GEN_2262; // @[util.scala 14:20:@5109.4]
  assign _T_1816 = $unsigned(_T_1815); // @[util.scala 14:20:@5110.4]
  assign _T_1817 = _T_1816[5:0]; // @[util.scala 14:20:@5111.4]
  assign _GEN_26 = _T_1817 % 6'h10; // @[util.scala 14:25:@5112.4]
  assign _T_1818 = _GEN_26[4:0]; // @[util.scala 14:25:@5112.4]
  assign _T_1819 = _T_1818 < _GEN_2263; // @[LoadQueue.scala 71:46:@5113.4]
  assign initBits_11 = _T_1819 & io_bbStart; // @[LoadQueue.scala 71:63:@5114.4]
  assign _T_1824 = 6'h1c - _GEN_2262; // @[util.scala 14:20:@5116.4]
  assign _T_1825 = $unsigned(_T_1824); // @[util.scala 14:20:@5117.4]
  assign _T_1826 = _T_1825[5:0]; // @[util.scala 14:20:@5118.4]
  assign _GEN_27 = _T_1826 % 6'h10; // @[util.scala 14:25:@5119.4]
  assign _T_1827 = _GEN_27[4:0]; // @[util.scala 14:25:@5119.4]
  assign _T_1828 = _T_1827 < _GEN_2263; // @[LoadQueue.scala 71:46:@5120.4]
  assign initBits_12 = _T_1828 & io_bbStart; // @[LoadQueue.scala 71:63:@5121.4]
  assign _T_1833 = 6'h1d - _GEN_2262; // @[util.scala 14:20:@5123.4]
  assign _T_1834 = $unsigned(_T_1833); // @[util.scala 14:20:@5124.4]
  assign _T_1835 = _T_1834[5:0]; // @[util.scala 14:20:@5125.4]
  assign _GEN_28 = _T_1835 % 6'h10; // @[util.scala 14:25:@5126.4]
  assign _T_1836 = _GEN_28[4:0]; // @[util.scala 14:25:@5126.4]
  assign _T_1837 = _T_1836 < _GEN_2263; // @[LoadQueue.scala 71:46:@5127.4]
  assign initBits_13 = _T_1837 & io_bbStart; // @[LoadQueue.scala 71:63:@5128.4]
  assign _T_1842 = 6'h1e - _GEN_2262; // @[util.scala 14:20:@5130.4]
  assign _T_1843 = $unsigned(_T_1842); // @[util.scala 14:20:@5131.4]
  assign _T_1844 = _T_1843[5:0]; // @[util.scala 14:20:@5132.4]
  assign _GEN_29 = _T_1844 % 6'h10; // @[util.scala 14:25:@5133.4]
  assign _T_1845 = _GEN_29[4:0]; // @[util.scala 14:25:@5133.4]
  assign _T_1846 = _T_1845 < _GEN_2263; // @[LoadQueue.scala 71:46:@5134.4]
  assign initBits_14 = _T_1846 & io_bbStart; // @[LoadQueue.scala 71:63:@5135.4]
  assign _T_1851 = 6'h1f - _GEN_2262; // @[util.scala 14:20:@5137.4]
  assign _T_1852 = $unsigned(_T_1851); // @[util.scala 14:20:@5138.4]
  assign _T_1853 = _T_1852[5:0]; // @[util.scala 14:20:@5139.4]
  assign _GEN_30 = _T_1853 % 6'h10; // @[util.scala 14:25:@5140.4]
  assign _T_1854 = _GEN_30[4:0]; // @[util.scala 14:25:@5140.4]
  assign _T_1855 = _T_1854 < _GEN_2263; // @[LoadQueue.scala 71:46:@5141.4]
  assign initBits_15 = _T_1855 & io_bbStart; // @[LoadQueue.scala 71:63:@5142.4]
  assign _T_1878 = allocatedEntries_0 | initBits_0; // @[LoadQueue.scala 73:78:@5160.4]
  assign _T_1879 = allocatedEntries_1 | initBits_1; // @[LoadQueue.scala 73:78:@5161.4]
  assign _T_1880 = allocatedEntries_2 | initBits_2; // @[LoadQueue.scala 73:78:@5162.4]
  assign _T_1881 = allocatedEntries_3 | initBits_3; // @[LoadQueue.scala 73:78:@5163.4]
  assign _T_1882 = allocatedEntries_4 | initBits_4; // @[LoadQueue.scala 73:78:@5164.4]
  assign _T_1883 = allocatedEntries_5 | initBits_5; // @[LoadQueue.scala 73:78:@5165.4]
  assign _T_1884 = allocatedEntries_6 | initBits_6; // @[LoadQueue.scala 73:78:@5166.4]
  assign _T_1885 = allocatedEntries_7 | initBits_7; // @[LoadQueue.scala 73:78:@5167.4]
  assign _T_1886 = allocatedEntries_8 | initBits_8; // @[LoadQueue.scala 73:78:@5168.4]
  assign _T_1887 = allocatedEntries_9 | initBits_9; // @[LoadQueue.scala 73:78:@5169.4]
  assign _T_1888 = allocatedEntries_10 | initBits_10; // @[LoadQueue.scala 73:78:@5170.4]
  assign _T_1889 = allocatedEntries_11 | initBits_11; // @[LoadQueue.scala 73:78:@5171.4]
  assign _T_1890 = allocatedEntries_12 | initBits_12; // @[LoadQueue.scala 73:78:@5172.4]
  assign _T_1891 = allocatedEntries_13 | initBits_13; // @[LoadQueue.scala 73:78:@5173.4]
  assign _T_1892 = allocatedEntries_14 | initBits_14; // @[LoadQueue.scala 73:78:@5174.4]
  assign _T_1893 = allocatedEntries_15 | initBits_15; // @[LoadQueue.scala 73:78:@5175.4]
  assign _T_1924 = _T_1719[3:0]; // @[:@5215.6]
  assign _GEN_1 = 4'h1 == _T_1924 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_2 = 4'h2 == _T_1924 ? io_bbLoadOffsets_2 : _GEN_1; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_3 = 4'h3 == _T_1924 ? io_bbLoadOffsets_3 : _GEN_2; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_4 = 4'h4 == _T_1924 ? io_bbLoadOffsets_4 : _GEN_3; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_5 = 4'h5 == _T_1924 ? io_bbLoadOffsets_5 : _GEN_4; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_6 = 4'h6 == _T_1924 ? io_bbLoadOffsets_6 : _GEN_5; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_7 = 4'h7 == _T_1924 ? io_bbLoadOffsets_7 : _GEN_6; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_8 = 4'h8 == _T_1924 ? io_bbLoadOffsets_8 : _GEN_7; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_9 = 4'h9 == _T_1924 ? io_bbLoadOffsets_9 : _GEN_8; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_10 = 4'ha == _T_1924 ? io_bbLoadOffsets_10 : _GEN_9; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_11 = 4'hb == _T_1924 ? io_bbLoadOffsets_11 : _GEN_10; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_12 = 4'hc == _T_1924 ? io_bbLoadOffsets_12 : _GEN_11; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_13 = 4'hd == _T_1924 ? io_bbLoadOffsets_13 : _GEN_12; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_14 = 4'he == _T_1924 ? io_bbLoadOffsets_14 : _GEN_13; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_15 = 4'hf == _T_1924 ? io_bbLoadOffsets_15 : _GEN_14; // @[LoadQueue.scala 77:20:@5216.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[LoadQueue.scala 76:25:@5209.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[LoadQueue.scala 76:25:@5209.4]
  assign _T_1942 = _T_1728[3:0]; // @[:@5231.6]
  assign _GEN_35 = 4'h1 == _T_1942 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_36 = 4'h2 == _T_1942 ? io_bbLoadOffsets_2 : _GEN_35; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_37 = 4'h3 == _T_1942 ? io_bbLoadOffsets_3 : _GEN_36; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_38 = 4'h4 == _T_1942 ? io_bbLoadOffsets_4 : _GEN_37; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_39 = 4'h5 == _T_1942 ? io_bbLoadOffsets_5 : _GEN_38; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_40 = 4'h6 == _T_1942 ? io_bbLoadOffsets_6 : _GEN_39; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_41 = 4'h7 == _T_1942 ? io_bbLoadOffsets_7 : _GEN_40; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_42 = 4'h8 == _T_1942 ? io_bbLoadOffsets_8 : _GEN_41; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_43 = 4'h9 == _T_1942 ? io_bbLoadOffsets_9 : _GEN_42; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_44 = 4'ha == _T_1942 ? io_bbLoadOffsets_10 : _GEN_43; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_45 = 4'hb == _T_1942 ? io_bbLoadOffsets_11 : _GEN_44; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_46 = 4'hc == _T_1942 ? io_bbLoadOffsets_12 : _GEN_45; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_47 = 4'hd == _T_1942 ? io_bbLoadOffsets_13 : _GEN_46; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_48 = 4'he == _T_1942 ? io_bbLoadOffsets_14 : _GEN_47; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_49 = 4'hf == _T_1942 ? io_bbLoadOffsets_15 : _GEN_48; // @[LoadQueue.scala 77:20:@5232.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[LoadQueue.scala 76:25:@5225.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[LoadQueue.scala 76:25:@5225.4]
  assign _T_1960 = _T_1737[3:0]; // @[:@5247.6]
  assign _GEN_69 = 4'h1 == _T_1960 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_70 = 4'h2 == _T_1960 ? io_bbLoadOffsets_2 : _GEN_69; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_71 = 4'h3 == _T_1960 ? io_bbLoadOffsets_3 : _GEN_70; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_72 = 4'h4 == _T_1960 ? io_bbLoadOffsets_4 : _GEN_71; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_73 = 4'h5 == _T_1960 ? io_bbLoadOffsets_5 : _GEN_72; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_74 = 4'h6 == _T_1960 ? io_bbLoadOffsets_6 : _GEN_73; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_75 = 4'h7 == _T_1960 ? io_bbLoadOffsets_7 : _GEN_74; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_76 = 4'h8 == _T_1960 ? io_bbLoadOffsets_8 : _GEN_75; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_77 = 4'h9 == _T_1960 ? io_bbLoadOffsets_9 : _GEN_76; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_78 = 4'ha == _T_1960 ? io_bbLoadOffsets_10 : _GEN_77; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_79 = 4'hb == _T_1960 ? io_bbLoadOffsets_11 : _GEN_78; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_80 = 4'hc == _T_1960 ? io_bbLoadOffsets_12 : _GEN_79; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_81 = 4'hd == _T_1960 ? io_bbLoadOffsets_13 : _GEN_80; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_82 = 4'he == _T_1960 ? io_bbLoadOffsets_14 : _GEN_81; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_83 = 4'hf == _T_1960 ? io_bbLoadOffsets_15 : _GEN_82; // @[LoadQueue.scala 77:20:@5248.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[LoadQueue.scala 76:25:@5241.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[LoadQueue.scala 76:25:@5241.4]
  assign _T_1978 = _T_1746[3:0]; // @[:@5263.6]
  assign _GEN_103 = 4'h1 == _T_1978 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_104 = 4'h2 == _T_1978 ? io_bbLoadOffsets_2 : _GEN_103; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_105 = 4'h3 == _T_1978 ? io_bbLoadOffsets_3 : _GEN_104; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_106 = 4'h4 == _T_1978 ? io_bbLoadOffsets_4 : _GEN_105; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_107 = 4'h5 == _T_1978 ? io_bbLoadOffsets_5 : _GEN_106; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_108 = 4'h6 == _T_1978 ? io_bbLoadOffsets_6 : _GEN_107; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_109 = 4'h7 == _T_1978 ? io_bbLoadOffsets_7 : _GEN_108; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_110 = 4'h8 == _T_1978 ? io_bbLoadOffsets_8 : _GEN_109; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_111 = 4'h9 == _T_1978 ? io_bbLoadOffsets_9 : _GEN_110; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_112 = 4'ha == _T_1978 ? io_bbLoadOffsets_10 : _GEN_111; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_113 = 4'hb == _T_1978 ? io_bbLoadOffsets_11 : _GEN_112; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_114 = 4'hc == _T_1978 ? io_bbLoadOffsets_12 : _GEN_113; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_115 = 4'hd == _T_1978 ? io_bbLoadOffsets_13 : _GEN_114; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_116 = 4'he == _T_1978 ? io_bbLoadOffsets_14 : _GEN_115; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_117 = 4'hf == _T_1978 ? io_bbLoadOffsets_15 : _GEN_116; // @[LoadQueue.scala 77:20:@5264.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[LoadQueue.scala 76:25:@5257.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[LoadQueue.scala 76:25:@5257.4]
  assign _T_1996 = _T_1755[3:0]; // @[:@5279.6]
  assign _GEN_137 = 4'h1 == _T_1996 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_138 = 4'h2 == _T_1996 ? io_bbLoadOffsets_2 : _GEN_137; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_139 = 4'h3 == _T_1996 ? io_bbLoadOffsets_3 : _GEN_138; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_140 = 4'h4 == _T_1996 ? io_bbLoadOffsets_4 : _GEN_139; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_141 = 4'h5 == _T_1996 ? io_bbLoadOffsets_5 : _GEN_140; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_142 = 4'h6 == _T_1996 ? io_bbLoadOffsets_6 : _GEN_141; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_143 = 4'h7 == _T_1996 ? io_bbLoadOffsets_7 : _GEN_142; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_144 = 4'h8 == _T_1996 ? io_bbLoadOffsets_8 : _GEN_143; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_145 = 4'h9 == _T_1996 ? io_bbLoadOffsets_9 : _GEN_144; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_146 = 4'ha == _T_1996 ? io_bbLoadOffsets_10 : _GEN_145; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_147 = 4'hb == _T_1996 ? io_bbLoadOffsets_11 : _GEN_146; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_148 = 4'hc == _T_1996 ? io_bbLoadOffsets_12 : _GEN_147; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_149 = 4'hd == _T_1996 ? io_bbLoadOffsets_13 : _GEN_148; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_150 = 4'he == _T_1996 ? io_bbLoadOffsets_14 : _GEN_149; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_151 = 4'hf == _T_1996 ? io_bbLoadOffsets_15 : _GEN_150; // @[LoadQueue.scala 77:20:@5280.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[LoadQueue.scala 76:25:@5273.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[LoadQueue.scala 76:25:@5273.4]
  assign _T_2014 = _T_1764[3:0]; // @[:@5295.6]
  assign _GEN_171 = 4'h1 == _T_2014 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_172 = 4'h2 == _T_2014 ? io_bbLoadOffsets_2 : _GEN_171; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_173 = 4'h3 == _T_2014 ? io_bbLoadOffsets_3 : _GEN_172; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_174 = 4'h4 == _T_2014 ? io_bbLoadOffsets_4 : _GEN_173; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_175 = 4'h5 == _T_2014 ? io_bbLoadOffsets_5 : _GEN_174; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_176 = 4'h6 == _T_2014 ? io_bbLoadOffsets_6 : _GEN_175; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_177 = 4'h7 == _T_2014 ? io_bbLoadOffsets_7 : _GEN_176; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_178 = 4'h8 == _T_2014 ? io_bbLoadOffsets_8 : _GEN_177; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_179 = 4'h9 == _T_2014 ? io_bbLoadOffsets_9 : _GEN_178; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_180 = 4'ha == _T_2014 ? io_bbLoadOffsets_10 : _GEN_179; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_181 = 4'hb == _T_2014 ? io_bbLoadOffsets_11 : _GEN_180; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_182 = 4'hc == _T_2014 ? io_bbLoadOffsets_12 : _GEN_181; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_183 = 4'hd == _T_2014 ? io_bbLoadOffsets_13 : _GEN_182; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_184 = 4'he == _T_2014 ? io_bbLoadOffsets_14 : _GEN_183; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_185 = 4'hf == _T_2014 ? io_bbLoadOffsets_15 : _GEN_184; // @[LoadQueue.scala 77:20:@5296.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[LoadQueue.scala 76:25:@5289.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[LoadQueue.scala 76:25:@5289.4]
  assign _T_2032 = _T_1773[3:0]; // @[:@5311.6]
  assign _GEN_205 = 4'h1 == _T_2032 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_206 = 4'h2 == _T_2032 ? io_bbLoadOffsets_2 : _GEN_205; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_207 = 4'h3 == _T_2032 ? io_bbLoadOffsets_3 : _GEN_206; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_208 = 4'h4 == _T_2032 ? io_bbLoadOffsets_4 : _GEN_207; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_209 = 4'h5 == _T_2032 ? io_bbLoadOffsets_5 : _GEN_208; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_210 = 4'h6 == _T_2032 ? io_bbLoadOffsets_6 : _GEN_209; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_211 = 4'h7 == _T_2032 ? io_bbLoadOffsets_7 : _GEN_210; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_212 = 4'h8 == _T_2032 ? io_bbLoadOffsets_8 : _GEN_211; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_213 = 4'h9 == _T_2032 ? io_bbLoadOffsets_9 : _GEN_212; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_214 = 4'ha == _T_2032 ? io_bbLoadOffsets_10 : _GEN_213; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_215 = 4'hb == _T_2032 ? io_bbLoadOffsets_11 : _GEN_214; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_216 = 4'hc == _T_2032 ? io_bbLoadOffsets_12 : _GEN_215; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_217 = 4'hd == _T_2032 ? io_bbLoadOffsets_13 : _GEN_216; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_218 = 4'he == _T_2032 ? io_bbLoadOffsets_14 : _GEN_217; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_219 = 4'hf == _T_2032 ? io_bbLoadOffsets_15 : _GEN_218; // @[LoadQueue.scala 77:20:@5312.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[LoadQueue.scala 76:25:@5305.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[LoadQueue.scala 76:25:@5305.4]
  assign _T_2050 = _T_1782[3:0]; // @[:@5327.6]
  assign _GEN_239 = 4'h1 == _T_2050 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_240 = 4'h2 == _T_2050 ? io_bbLoadOffsets_2 : _GEN_239; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_241 = 4'h3 == _T_2050 ? io_bbLoadOffsets_3 : _GEN_240; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_242 = 4'h4 == _T_2050 ? io_bbLoadOffsets_4 : _GEN_241; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_243 = 4'h5 == _T_2050 ? io_bbLoadOffsets_5 : _GEN_242; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_244 = 4'h6 == _T_2050 ? io_bbLoadOffsets_6 : _GEN_243; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_245 = 4'h7 == _T_2050 ? io_bbLoadOffsets_7 : _GEN_244; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_246 = 4'h8 == _T_2050 ? io_bbLoadOffsets_8 : _GEN_245; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_247 = 4'h9 == _T_2050 ? io_bbLoadOffsets_9 : _GEN_246; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_248 = 4'ha == _T_2050 ? io_bbLoadOffsets_10 : _GEN_247; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_249 = 4'hb == _T_2050 ? io_bbLoadOffsets_11 : _GEN_248; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_250 = 4'hc == _T_2050 ? io_bbLoadOffsets_12 : _GEN_249; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_251 = 4'hd == _T_2050 ? io_bbLoadOffsets_13 : _GEN_250; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_252 = 4'he == _T_2050 ? io_bbLoadOffsets_14 : _GEN_251; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_253 = 4'hf == _T_2050 ? io_bbLoadOffsets_15 : _GEN_252; // @[LoadQueue.scala 77:20:@5328.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[LoadQueue.scala 76:25:@5321.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[LoadQueue.scala 76:25:@5321.4]
  assign _T_2068 = _T_1791[3:0]; // @[:@5343.6]
  assign _GEN_273 = 4'h1 == _T_2068 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_274 = 4'h2 == _T_2068 ? io_bbLoadOffsets_2 : _GEN_273; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_275 = 4'h3 == _T_2068 ? io_bbLoadOffsets_3 : _GEN_274; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_276 = 4'h4 == _T_2068 ? io_bbLoadOffsets_4 : _GEN_275; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_277 = 4'h5 == _T_2068 ? io_bbLoadOffsets_5 : _GEN_276; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_278 = 4'h6 == _T_2068 ? io_bbLoadOffsets_6 : _GEN_277; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_279 = 4'h7 == _T_2068 ? io_bbLoadOffsets_7 : _GEN_278; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_280 = 4'h8 == _T_2068 ? io_bbLoadOffsets_8 : _GEN_279; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_281 = 4'h9 == _T_2068 ? io_bbLoadOffsets_9 : _GEN_280; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_282 = 4'ha == _T_2068 ? io_bbLoadOffsets_10 : _GEN_281; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_283 = 4'hb == _T_2068 ? io_bbLoadOffsets_11 : _GEN_282; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_284 = 4'hc == _T_2068 ? io_bbLoadOffsets_12 : _GEN_283; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_285 = 4'hd == _T_2068 ? io_bbLoadOffsets_13 : _GEN_284; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_286 = 4'he == _T_2068 ? io_bbLoadOffsets_14 : _GEN_285; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_287 = 4'hf == _T_2068 ? io_bbLoadOffsets_15 : _GEN_286; // @[LoadQueue.scala 77:20:@5344.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[LoadQueue.scala 76:25:@5337.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[LoadQueue.scala 76:25:@5337.4]
  assign _T_2086 = _T_1800[3:0]; // @[:@5359.6]
  assign _GEN_307 = 4'h1 == _T_2086 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_308 = 4'h2 == _T_2086 ? io_bbLoadOffsets_2 : _GEN_307; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_309 = 4'h3 == _T_2086 ? io_bbLoadOffsets_3 : _GEN_308; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_310 = 4'h4 == _T_2086 ? io_bbLoadOffsets_4 : _GEN_309; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_311 = 4'h5 == _T_2086 ? io_bbLoadOffsets_5 : _GEN_310; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_312 = 4'h6 == _T_2086 ? io_bbLoadOffsets_6 : _GEN_311; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_313 = 4'h7 == _T_2086 ? io_bbLoadOffsets_7 : _GEN_312; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_314 = 4'h8 == _T_2086 ? io_bbLoadOffsets_8 : _GEN_313; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_315 = 4'h9 == _T_2086 ? io_bbLoadOffsets_9 : _GEN_314; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_316 = 4'ha == _T_2086 ? io_bbLoadOffsets_10 : _GEN_315; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_317 = 4'hb == _T_2086 ? io_bbLoadOffsets_11 : _GEN_316; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_318 = 4'hc == _T_2086 ? io_bbLoadOffsets_12 : _GEN_317; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_319 = 4'hd == _T_2086 ? io_bbLoadOffsets_13 : _GEN_318; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_320 = 4'he == _T_2086 ? io_bbLoadOffsets_14 : _GEN_319; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_321 = 4'hf == _T_2086 ? io_bbLoadOffsets_15 : _GEN_320; // @[LoadQueue.scala 77:20:@5360.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[LoadQueue.scala 76:25:@5353.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[LoadQueue.scala 76:25:@5353.4]
  assign _T_2104 = _T_1809[3:0]; // @[:@5375.6]
  assign _GEN_341 = 4'h1 == _T_2104 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_342 = 4'h2 == _T_2104 ? io_bbLoadOffsets_2 : _GEN_341; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_343 = 4'h3 == _T_2104 ? io_bbLoadOffsets_3 : _GEN_342; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_344 = 4'h4 == _T_2104 ? io_bbLoadOffsets_4 : _GEN_343; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_345 = 4'h5 == _T_2104 ? io_bbLoadOffsets_5 : _GEN_344; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_346 = 4'h6 == _T_2104 ? io_bbLoadOffsets_6 : _GEN_345; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_347 = 4'h7 == _T_2104 ? io_bbLoadOffsets_7 : _GEN_346; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_348 = 4'h8 == _T_2104 ? io_bbLoadOffsets_8 : _GEN_347; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_349 = 4'h9 == _T_2104 ? io_bbLoadOffsets_9 : _GEN_348; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_350 = 4'ha == _T_2104 ? io_bbLoadOffsets_10 : _GEN_349; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_351 = 4'hb == _T_2104 ? io_bbLoadOffsets_11 : _GEN_350; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_352 = 4'hc == _T_2104 ? io_bbLoadOffsets_12 : _GEN_351; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_353 = 4'hd == _T_2104 ? io_bbLoadOffsets_13 : _GEN_352; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_354 = 4'he == _T_2104 ? io_bbLoadOffsets_14 : _GEN_353; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_355 = 4'hf == _T_2104 ? io_bbLoadOffsets_15 : _GEN_354; // @[LoadQueue.scala 77:20:@5376.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[LoadQueue.scala 76:25:@5369.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[LoadQueue.scala 76:25:@5369.4]
  assign _T_2122 = _T_1818[3:0]; // @[:@5391.6]
  assign _GEN_375 = 4'h1 == _T_2122 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_376 = 4'h2 == _T_2122 ? io_bbLoadOffsets_2 : _GEN_375; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_377 = 4'h3 == _T_2122 ? io_bbLoadOffsets_3 : _GEN_376; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_378 = 4'h4 == _T_2122 ? io_bbLoadOffsets_4 : _GEN_377; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_379 = 4'h5 == _T_2122 ? io_bbLoadOffsets_5 : _GEN_378; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_380 = 4'h6 == _T_2122 ? io_bbLoadOffsets_6 : _GEN_379; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_381 = 4'h7 == _T_2122 ? io_bbLoadOffsets_7 : _GEN_380; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_382 = 4'h8 == _T_2122 ? io_bbLoadOffsets_8 : _GEN_381; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_383 = 4'h9 == _T_2122 ? io_bbLoadOffsets_9 : _GEN_382; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_384 = 4'ha == _T_2122 ? io_bbLoadOffsets_10 : _GEN_383; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_385 = 4'hb == _T_2122 ? io_bbLoadOffsets_11 : _GEN_384; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_386 = 4'hc == _T_2122 ? io_bbLoadOffsets_12 : _GEN_385; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_387 = 4'hd == _T_2122 ? io_bbLoadOffsets_13 : _GEN_386; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_388 = 4'he == _T_2122 ? io_bbLoadOffsets_14 : _GEN_387; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_389 = 4'hf == _T_2122 ? io_bbLoadOffsets_15 : _GEN_388; // @[LoadQueue.scala 77:20:@5392.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[LoadQueue.scala 76:25:@5385.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[LoadQueue.scala 76:25:@5385.4]
  assign _T_2140 = _T_1827[3:0]; // @[:@5407.6]
  assign _GEN_409 = 4'h1 == _T_2140 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_410 = 4'h2 == _T_2140 ? io_bbLoadOffsets_2 : _GEN_409; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_411 = 4'h3 == _T_2140 ? io_bbLoadOffsets_3 : _GEN_410; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_412 = 4'h4 == _T_2140 ? io_bbLoadOffsets_4 : _GEN_411; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_413 = 4'h5 == _T_2140 ? io_bbLoadOffsets_5 : _GEN_412; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_414 = 4'h6 == _T_2140 ? io_bbLoadOffsets_6 : _GEN_413; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_415 = 4'h7 == _T_2140 ? io_bbLoadOffsets_7 : _GEN_414; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_416 = 4'h8 == _T_2140 ? io_bbLoadOffsets_8 : _GEN_415; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_417 = 4'h9 == _T_2140 ? io_bbLoadOffsets_9 : _GEN_416; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_418 = 4'ha == _T_2140 ? io_bbLoadOffsets_10 : _GEN_417; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_419 = 4'hb == _T_2140 ? io_bbLoadOffsets_11 : _GEN_418; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_420 = 4'hc == _T_2140 ? io_bbLoadOffsets_12 : _GEN_419; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_421 = 4'hd == _T_2140 ? io_bbLoadOffsets_13 : _GEN_420; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_422 = 4'he == _T_2140 ? io_bbLoadOffsets_14 : _GEN_421; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_423 = 4'hf == _T_2140 ? io_bbLoadOffsets_15 : _GEN_422; // @[LoadQueue.scala 77:20:@5408.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[LoadQueue.scala 76:25:@5401.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[LoadQueue.scala 76:25:@5401.4]
  assign _T_2158 = _T_1836[3:0]; // @[:@5423.6]
  assign _GEN_443 = 4'h1 == _T_2158 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_444 = 4'h2 == _T_2158 ? io_bbLoadOffsets_2 : _GEN_443; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_445 = 4'h3 == _T_2158 ? io_bbLoadOffsets_3 : _GEN_444; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_446 = 4'h4 == _T_2158 ? io_bbLoadOffsets_4 : _GEN_445; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_447 = 4'h5 == _T_2158 ? io_bbLoadOffsets_5 : _GEN_446; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_448 = 4'h6 == _T_2158 ? io_bbLoadOffsets_6 : _GEN_447; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_449 = 4'h7 == _T_2158 ? io_bbLoadOffsets_7 : _GEN_448; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_450 = 4'h8 == _T_2158 ? io_bbLoadOffsets_8 : _GEN_449; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_451 = 4'h9 == _T_2158 ? io_bbLoadOffsets_9 : _GEN_450; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_452 = 4'ha == _T_2158 ? io_bbLoadOffsets_10 : _GEN_451; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_453 = 4'hb == _T_2158 ? io_bbLoadOffsets_11 : _GEN_452; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_454 = 4'hc == _T_2158 ? io_bbLoadOffsets_12 : _GEN_453; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_455 = 4'hd == _T_2158 ? io_bbLoadOffsets_13 : _GEN_454; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_456 = 4'he == _T_2158 ? io_bbLoadOffsets_14 : _GEN_455; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_457 = 4'hf == _T_2158 ? io_bbLoadOffsets_15 : _GEN_456; // @[LoadQueue.scala 77:20:@5424.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[LoadQueue.scala 76:25:@5417.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[LoadQueue.scala 76:25:@5417.4]
  assign _T_2176 = _T_1845[3:0]; // @[:@5439.6]
  assign _GEN_477 = 4'h1 == _T_2176 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_478 = 4'h2 == _T_2176 ? io_bbLoadOffsets_2 : _GEN_477; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_479 = 4'h3 == _T_2176 ? io_bbLoadOffsets_3 : _GEN_478; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_480 = 4'h4 == _T_2176 ? io_bbLoadOffsets_4 : _GEN_479; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_481 = 4'h5 == _T_2176 ? io_bbLoadOffsets_5 : _GEN_480; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_482 = 4'h6 == _T_2176 ? io_bbLoadOffsets_6 : _GEN_481; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_483 = 4'h7 == _T_2176 ? io_bbLoadOffsets_7 : _GEN_482; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_484 = 4'h8 == _T_2176 ? io_bbLoadOffsets_8 : _GEN_483; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_485 = 4'h9 == _T_2176 ? io_bbLoadOffsets_9 : _GEN_484; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_486 = 4'ha == _T_2176 ? io_bbLoadOffsets_10 : _GEN_485; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_487 = 4'hb == _T_2176 ? io_bbLoadOffsets_11 : _GEN_486; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_488 = 4'hc == _T_2176 ? io_bbLoadOffsets_12 : _GEN_487; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_489 = 4'hd == _T_2176 ? io_bbLoadOffsets_13 : _GEN_488; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_490 = 4'he == _T_2176 ? io_bbLoadOffsets_14 : _GEN_489; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_491 = 4'hf == _T_2176 ? io_bbLoadOffsets_15 : _GEN_490; // @[LoadQueue.scala 77:20:@5440.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[LoadQueue.scala 76:25:@5433.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[LoadQueue.scala 76:25:@5433.4]
  assign _T_2194 = _T_1854[3:0]; // @[:@5455.6]
  assign _GEN_511 = 4'h1 == _T_2194 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_512 = 4'h2 == _T_2194 ? io_bbLoadOffsets_2 : _GEN_511; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_513 = 4'h3 == _T_2194 ? io_bbLoadOffsets_3 : _GEN_512; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_514 = 4'h4 == _T_2194 ? io_bbLoadOffsets_4 : _GEN_513; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_515 = 4'h5 == _T_2194 ? io_bbLoadOffsets_5 : _GEN_514; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_516 = 4'h6 == _T_2194 ? io_bbLoadOffsets_6 : _GEN_515; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_517 = 4'h7 == _T_2194 ? io_bbLoadOffsets_7 : _GEN_516; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_518 = 4'h8 == _T_2194 ? io_bbLoadOffsets_8 : _GEN_517; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_519 = 4'h9 == _T_2194 ? io_bbLoadOffsets_9 : _GEN_518; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_520 = 4'ha == _T_2194 ? io_bbLoadOffsets_10 : _GEN_519; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_521 = 4'hb == _T_2194 ? io_bbLoadOffsets_11 : _GEN_520; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_522 = 4'hc == _T_2194 ? io_bbLoadOffsets_12 : _GEN_521; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_523 = 4'hd == _T_2194 ? io_bbLoadOffsets_13 : _GEN_522; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_524 = 4'he == _T_2194 ? io_bbLoadOffsets_14 : _GEN_523; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_525 = 4'hf == _T_2194 ? io_bbLoadOffsets_15 : _GEN_524; // @[LoadQueue.scala 77:20:@5456.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[LoadQueue.scala 76:25:@5449.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[LoadQueue.scala 76:25:@5449.4]
  assign _T_2216 = _GEN_15 + 4'h1; // @[util.scala 10:8:@5474.6]
  assign _GEN_31 = _T_2216 % 5'h10; // @[util.scala 10:14:@5475.6]
  assign _T_2217 = _GEN_31[4:0]; // @[util.scala 10:14:@5475.6]
  assign _GEN_2327 = {{1'd0}, io_storeTail}; // @[LoadQueue.scala 97:56:@5476.6]
  assign _T_2218 = _T_2217 == _GEN_2327; // @[LoadQueue.scala 97:56:@5476.6]
  assign _T_2219 = io_storeEmpty & _T_2218; // @[LoadQueue.scala 96:50:@5477.6]
  assign _T_2221 = _T_2219 == 1'h0; // @[LoadQueue.scala 96:34:@5478.6]
  assign _T_2223 = previousStoreHead <= offsetQ_0; // @[LoadQueue.scala 101:36:@5486.8]
  assign _T_2224 = offsetQ_0 < io_storeHead; // @[LoadQueue.scala 101:86:@5487.8]
  assign _T_2225 = _T_2223 & _T_2224; // @[LoadQueue.scala 101:61:@5488.8]
  assign _T_2227 = previousStoreHead > io_storeHead; // @[LoadQueue.scala 103:36:@5493.10]
  assign _T_2228 = io_storeHead <= offsetQ_0; // @[LoadQueue.scala 103:69:@5494.10]
  assign _T_2229 = offsetQ_0 < previousStoreHead; // @[LoadQueue.scala 104:31:@5495.10]
  assign _T_2230 = _T_2228 & _T_2229; // @[LoadQueue.scala 103:94:@5496.10]
  assign _T_2232 = _T_2230 == 1'h0; // @[LoadQueue.scala 103:54:@5497.10]
  assign _T_2233 = _T_2227 & _T_2232; // @[LoadQueue.scala 103:51:@5498.10]
  assign _GEN_560 = _T_2233 ? 1'h0 : checkBits_0; // @[LoadQueue.scala 104:53:@5499.10]
  assign _GEN_561 = _T_2225 ? 1'h0 : _GEN_560; // @[LoadQueue.scala 101:102:@5489.8]
  assign _GEN_562 = io_storeEmpty ? 1'h0 : _GEN_561; // @[LoadQueue.scala 99:27:@5482.6]
  assign _GEN_563 = initBits_0 ? _T_2221 : _GEN_562; // @[LoadQueue.scala 95:34:@5467.4]
  assign _T_2246 = _GEN_49 + 4'h1; // @[util.scala 10:8:@5510.6]
  assign _GEN_34 = _T_2246 % 5'h10; // @[util.scala 10:14:@5511.6]
  assign _T_2247 = _GEN_34[4:0]; // @[util.scala 10:14:@5511.6]
  assign _T_2248 = _T_2247 == _GEN_2327; // @[LoadQueue.scala 97:56:@5512.6]
  assign _T_2249 = io_storeEmpty & _T_2248; // @[LoadQueue.scala 96:50:@5513.6]
  assign _T_2251 = _T_2249 == 1'h0; // @[LoadQueue.scala 96:34:@5514.6]
  assign _T_2253 = previousStoreHead <= offsetQ_1; // @[LoadQueue.scala 101:36:@5522.8]
  assign _T_2254 = offsetQ_1 < io_storeHead; // @[LoadQueue.scala 101:86:@5523.8]
  assign _T_2255 = _T_2253 & _T_2254; // @[LoadQueue.scala 101:61:@5524.8]
  assign _T_2258 = io_storeHead <= offsetQ_1; // @[LoadQueue.scala 103:69:@5530.10]
  assign _T_2259 = offsetQ_1 < previousStoreHead; // @[LoadQueue.scala 104:31:@5531.10]
  assign _T_2260 = _T_2258 & _T_2259; // @[LoadQueue.scala 103:94:@5532.10]
  assign _T_2262 = _T_2260 == 1'h0; // @[LoadQueue.scala 103:54:@5533.10]
  assign _T_2263 = _T_2227 & _T_2262; // @[LoadQueue.scala 103:51:@5534.10]
  assign _GEN_580 = _T_2263 ? 1'h0 : checkBits_1; // @[LoadQueue.scala 104:53:@5535.10]
  assign _GEN_581 = _T_2255 ? 1'h0 : _GEN_580; // @[LoadQueue.scala 101:102:@5525.8]
  assign _GEN_582 = io_storeEmpty ? 1'h0 : _GEN_581; // @[LoadQueue.scala 99:27:@5518.6]
  assign _GEN_583 = initBits_1 ? _T_2251 : _GEN_582; // @[LoadQueue.scala 95:34:@5503.4]
  assign _T_2276 = _GEN_83 + 4'h1; // @[util.scala 10:8:@5546.6]
  assign _GEN_50 = _T_2276 % 5'h10; // @[util.scala 10:14:@5547.6]
  assign _T_2277 = _GEN_50[4:0]; // @[util.scala 10:14:@5547.6]
  assign _T_2278 = _T_2277 == _GEN_2327; // @[LoadQueue.scala 97:56:@5548.6]
  assign _T_2279 = io_storeEmpty & _T_2278; // @[LoadQueue.scala 96:50:@5549.6]
  assign _T_2281 = _T_2279 == 1'h0; // @[LoadQueue.scala 96:34:@5550.6]
  assign _T_2283 = previousStoreHead <= offsetQ_2; // @[LoadQueue.scala 101:36:@5558.8]
  assign _T_2284 = offsetQ_2 < io_storeHead; // @[LoadQueue.scala 101:86:@5559.8]
  assign _T_2285 = _T_2283 & _T_2284; // @[LoadQueue.scala 101:61:@5560.8]
  assign _T_2288 = io_storeHead <= offsetQ_2; // @[LoadQueue.scala 103:69:@5566.10]
  assign _T_2289 = offsetQ_2 < previousStoreHead; // @[LoadQueue.scala 104:31:@5567.10]
  assign _T_2290 = _T_2288 & _T_2289; // @[LoadQueue.scala 103:94:@5568.10]
  assign _T_2292 = _T_2290 == 1'h0; // @[LoadQueue.scala 103:54:@5569.10]
  assign _T_2293 = _T_2227 & _T_2292; // @[LoadQueue.scala 103:51:@5570.10]
  assign _GEN_600 = _T_2293 ? 1'h0 : checkBits_2; // @[LoadQueue.scala 104:53:@5571.10]
  assign _GEN_601 = _T_2285 ? 1'h0 : _GEN_600; // @[LoadQueue.scala 101:102:@5561.8]
  assign _GEN_602 = io_storeEmpty ? 1'h0 : _GEN_601; // @[LoadQueue.scala 99:27:@5554.6]
  assign _GEN_603 = initBits_2 ? _T_2281 : _GEN_602; // @[LoadQueue.scala 95:34:@5539.4]
  assign _T_2306 = _GEN_117 + 4'h1; // @[util.scala 10:8:@5582.6]
  assign _GEN_51 = _T_2306 % 5'h10; // @[util.scala 10:14:@5583.6]
  assign _T_2307 = _GEN_51[4:0]; // @[util.scala 10:14:@5583.6]
  assign _T_2308 = _T_2307 == _GEN_2327; // @[LoadQueue.scala 97:56:@5584.6]
  assign _T_2309 = io_storeEmpty & _T_2308; // @[LoadQueue.scala 96:50:@5585.6]
  assign _T_2311 = _T_2309 == 1'h0; // @[LoadQueue.scala 96:34:@5586.6]
  assign _T_2313 = previousStoreHead <= offsetQ_3; // @[LoadQueue.scala 101:36:@5594.8]
  assign _T_2314 = offsetQ_3 < io_storeHead; // @[LoadQueue.scala 101:86:@5595.8]
  assign _T_2315 = _T_2313 & _T_2314; // @[LoadQueue.scala 101:61:@5596.8]
  assign _T_2318 = io_storeHead <= offsetQ_3; // @[LoadQueue.scala 103:69:@5602.10]
  assign _T_2319 = offsetQ_3 < previousStoreHead; // @[LoadQueue.scala 104:31:@5603.10]
  assign _T_2320 = _T_2318 & _T_2319; // @[LoadQueue.scala 103:94:@5604.10]
  assign _T_2322 = _T_2320 == 1'h0; // @[LoadQueue.scala 103:54:@5605.10]
  assign _T_2323 = _T_2227 & _T_2322; // @[LoadQueue.scala 103:51:@5606.10]
  assign _GEN_620 = _T_2323 ? 1'h0 : checkBits_3; // @[LoadQueue.scala 104:53:@5607.10]
  assign _GEN_621 = _T_2315 ? 1'h0 : _GEN_620; // @[LoadQueue.scala 101:102:@5597.8]
  assign _GEN_622 = io_storeEmpty ? 1'h0 : _GEN_621; // @[LoadQueue.scala 99:27:@5590.6]
  assign _GEN_623 = initBits_3 ? _T_2311 : _GEN_622; // @[LoadQueue.scala 95:34:@5575.4]
  assign _T_2336 = _GEN_151 + 4'h1; // @[util.scala 10:8:@5618.6]
  assign _GEN_52 = _T_2336 % 5'h10; // @[util.scala 10:14:@5619.6]
  assign _T_2337 = _GEN_52[4:0]; // @[util.scala 10:14:@5619.6]
  assign _T_2338 = _T_2337 == _GEN_2327; // @[LoadQueue.scala 97:56:@5620.6]
  assign _T_2339 = io_storeEmpty & _T_2338; // @[LoadQueue.scala 96:50:@5621.6]
  assign _T_2341 = _T_2339 == 1'h0; // @[LoadQueue.scala 96:34:@5622.6]
  assign _T_2343 = previousStoreHead <= offsetQ_4; // @[LoadQueue.scala 101:36:@5630.8]
  assign _T_2344 = offsetQ_4 < io_storeHead; // @[LoadQueue.scala 101:86:@5631.8]
  assign _T_2345 = _T_2343 & _T_2344; // @[LoadQueue.scala 101:61:@5632.8]
  assign _T_2348 = io_storeHead <= offsetQ_4; // @[LoadQueue.scala 103:69:@5638.10]
  assign _T_2349 = offsetQ_4 < previousStoreHead; // @[LoadQueue.scala 104:31:@5639.10]
  assign _T_2350 = _T_2348 & _T_2349; // @[LoadQueue.scala 103:94:@5640.10]
  assign _T_2352 = _T_2350 == 1'h0; // @[LoadQueue.scala 103:54:@5641.10]
  assign _T_2353 = _T_2227 & _T_2352; // @[LoadQueue.scala 103:51:@5642.10]
  assign _GEN_640 = _T_2353 ? 1'h0 : checkBits_4; // @[LoadQueue.scala 104:53:@5643.10]
  assign _GEN_641 = _T_2345 ? 1'h0 : _GEN_640; // @[LoadQueue.scala 101:102:@5633.8]
  assign _GEN_642 = io_storeEmpty ? 1'h0 : _GEN_641; // @[LoadQueue.scala 99:27:@5626.6]
  assign _GEN_643 = initBits_4 ? _T_2341 : _GEN_642; // @[LoadQueue.scala 95:34:@5611.4]
  assign _T_2366 = _GEN_185 + 4'h1; // @[util.scala 10:8:@5654.6]
  assign _GEN_53 = _T_2366 % 5'h10; // @[util.scala 10:14:@5655.6]
  assign _T_2367 = _GEN_53[4:0]; // @[util.scala 10:14:@5655.6]
  assign _T_2368 = _T_2367 == _GEN_2327; // @[LoadQueue.scala 97:56:@5656.6]
  assign _T_2369 = io_storeEmpty & _T_2368; // @[LoadQueue.scala 96:50:@5657.6]
  assign _T_2371 = _T_2369 == 1'h0; // @[LoadQueue.scala 96:34:@5658.6]
  assign _T_2373 = previousStoreHead <= offsetQ_5; // @[LoadQueue.scala 101:36:@5666.8]
  assign _T_2374 = offsetQ_5 < io_storeHead; // @[LoadQueue.scala 101:86:@5667.8]
  assign _T_2375 = _T_2373 & _T_2374; // @[LoadQueue.scala 101:61:@5668.8]
  assign _T_2378 = io_storeHead <= offsetQ_5; // @[LoadQueue.scala 103:69:@5674.10]
  assign _T_2379 = offsetQ_5 < previousStoreHead; // @[LoadQueue.scala 104:31:@5675.10]
  assign _T_2380 = _T_2378 & _T_2379; // @[LoadQueue.scala 103:94:@5676.10]
  assign _T_2382 = _T_2380 == 1'h0; // @[LoadQueue.scala 103:54:@5677.10]
  assign _T_2383 = _T_2227 & _T_2382; // @[LoadQueue.scala 103:51:@5678.10]
  assign _GEN_660 = _T_2383 ? 1'h0 : checkBits_5; // @[LoadQueue.scala 104:53:@5679.10]
  assign _GEN_661 = _T_2375 ? 1'h0 : _GEN_660; // @[LoadQueue.scala 101:102:@5669.8]
  assign _GEN_662 = io_storeEmpty ? 1'h0 : _GEN_661; // @[LoadQueue.scala 99:27:@5662.6]
  assign _GEN_663 = initBits_5 ? _T_2371 : _GEN_662; // @[LoadQueue.scala 95:34:@5647.4]
  assign _T_2396 = _GEN_219 + 4'h1; // @[util.scala 10:8:@5690.6]
  assign _GEN_54 = _T_2396 % 5'h10; // @[util.scala 10:14:@5691.6]
  assign _T_2397 = _GEN_54[4:0]; // @[util.scala 10:14:@5691.6]
  assign _T_2398 = _T_2397 == _GEN_2327; // @[LoadQueue.scala 97:56:@5692.6]
  assign _T_2399 = io_storeEmpty & _T_2398; // @[LoadQueue.scala 96:50:@5693.6]
  assign _T_2401 = _T_2399 == 1'h0; // @[LoadQueue.scala 96:34:@5694.6]
  assign _T_2403 = previousStoreHead <= offsetQ_6; // @[LoadQueue.scala 101:36:@5702.8]
  assign _T_2404 = offsetQ_6 < io_storeHead; // @[LoadQueue.scala 101:86:@5703.8]
  assign _T_2405 = _T_2403 & _T_2404; // @[LoadQueue.scala 101:61:@5704.8]
  assign _T_2408 = io_storeHead <= offsetQ_6; // @[LoadQueue.scala 103:69:@5710.10]
  assign _T_2409 = offsetQ_6 < previousStoreHead; // @[LoadQueue.scala 104:31:@5711.10]
  assign _T_2410 = _T_2408 & _T_2409; // @[LoadQueue.scala 103:94:@5712.10]
  assign _T_2412 = _T_2410 == 1'h0; // @[LoadQueue.scala 103:54:@5713.10]
  assign _T_2413 = _T_2227 & _T_2412; // @[LoadQueue.scala 103:51:@5714.10]
  assign _GEN_680 = _T_2413 ? 1'h0 : checkBits_6; // @[LoadQueue.scala 104:53:@5715.10]
  assign _GEN_681 = _T_2405 ? 1'h0 : _GEN_680; // @[LoadQueue.scala 101:102:@5705.8]
  assign _GEN_682 = io_storeEmpty ? 1'h0 : _GEN_681; // @[LoadQueue.scala 99:27:@5698.6]
  assign _GEN_683 = initBits_6 ? _T_2401 : _GEN_682; // @[LoadQueue.scala 95:34:@5683.4]
  assign _T_2426 = _GEN_253 + 4'h1; // @[util.scala 10:8:@5726.6]
  assign _GEN_55 = _T_2426 % 5'h10; // @[util.scala 10:14:@5727.6]
  assign _T_2427 = _GEN_55[4:0]; // @[util.scala 10:14:@5727.6]
  assign _T_2428 = _T_2427 == _GEN_2327; // @[LoadQueue.scala 97:56:@5728.6]
  assign _T_2429 = io_storeEmpty & _T_2428; // @[LoadQueue.scala 96:50:@5729.6]
  assign _T_2431 = _T_2429 == 1'h0; // @[LoadQueue.scala 96:34:@5730.6]
  assign _T_2433 = previousStoreHead <= offsetQ_7; // @[LoadQueue.scala 101:36:@5738.8]
  assign _T_2434 = offsetQ_7 < io_storeHead; // @[LoadQueue.scala 101:86:@5739.8]
  assign _T_2435 = _T_2433 & _T_2434; // @[LoadQueue.scala 101:61:@5740.8]
  assign _T_2438 = io_storeHead <= offsetQ_7; // @[LoadQueue.scala 103:69:@5746.10]
  assign _T_2439 = offsetQ_7 < previousStoreHead; // @[LoadQueue.scala 104:31:@5747.10]
  assign _T_2440 = _T_2438 & _T_2439; // @[LoadQueue.scala 103:94:@5748.10]
  assign _T_2442 = _T_2440 == 1'h0; // @[LoadQueue.scala 103:54:@5749.10]
  assign _T_2443 = _T_2227 & _T_2442; // @[LoadQueue.scala 103:51:@5750.10]
  assign _GEN_700 = _T_2443 ? 1'h0 : checkBits_7; // @[LoadQueue.scala 104:53:@5751.10]
  assign _GEN_701 = _T_2435 ? 1'h0 : _GEN_700; // @[LoadQueue.scala 101:102:@5741.8]
  assign _GEN_702 = io_storeEmpty ? 1'h0 : _GEN_701; // @[LoadQueue.scala 99:27:@5734.6]
  assign _GEN_703 = initBits_7 ? _T_2431 : _GEN_702; // @[LoadQueue.scala 95:34:@5719.4]
  assign _T_2456 = _GEN_287 + 4'h1; // @[util.scala 10:8:@5762.6]
  assign _GEN_56 = _T_2456 % 5'h10; // @[util.scala 10:14:@5763.6]
  assign _T_2457 = _GEN_56[4:0]; // @[util.scala 10:14:@5763.6]
  assign _T_2458 = _T_2457 == _GEN_2327; // @[LoadQueue.scala 97:56:@5764.6]
  assign _T_2459 = io_storeEmpty & _T_2458; // @[LoadQueue.scala 96:50:@5765.6]
  assign _T_2461 = _T_2459 == 1'h0; // @[LoadQueue.scala 96:34:@5766.6]
  assign _T_2463 = previousStoreHead <= offsetQ_8; // @[LoadQueue.scala 101:36:@5774.8]
  assign _T_2464 = offsetQ_8 < io_storeHead; // @[LoadQueue.scala 101:86:@5775.8]
  assign _T_2465 = _T_2463 & _T_2464; // @[LoadQueue.scala 101:61:@5776.8]
  assign _T_2468 = io_storeHead <= offsetQ_8; // @[LoadQueue.scala 103:69:@5782.10]
  assign _T_2469 = offsetQ_8 < previousStoreHead; // @[LoadQueue.scala 104:31:@5783.10]
  assign _T_2470 = _T_2468 & _T_2469; // @[LoadQueue.scala 103:94:@5784.10]
  assign _T_2472 = _T_2470 == 1'h0; // @[LoadQueue.scala 103:54:@5785.10]
  assign _T_2473 = _T_2227 & _T_2472; // @[LoadQueue.scala 103:51:@5786.10]
  assign _GEN_720 = _T_2473 ? 1'h0 : checkBits_8; // @[LoadQueue.scala 104:53:@5787.10]
  assign _GEN_721 = _T_2465 ? 1'h0 : _GEN_720; // @[LoadQueue.scala 101:102:@5777.8]
  assign _GEN_722 = io_storeEmpty ? 1'h0 : _GEN_721; // @[LoadQueue.scala 99:27:@5770.6]
  assign _GEN_723 = initBits_8 ? _T_2461 : _GEN_722; // @[LoadQueue.scala 95:34:@5755.4]
  assign _T_2486 = _GEN_321 + 4'h1; // @[util.scala 10:8:@5798.6]
  assign _GEN_57 = _T_2486 % 5'h10; // @[util.scala 10:14:@5799.6]
  assign _T_2487 = _GEN_57[4:0]; // @[util.scala 10:14:@5799.6]
  assign _T_2488 = _T_2487 == _GEN_2327; // @[LoadQueue.scala 97:56:@5800.6]
  assign _T_2489 = io_storeEmpty & _T_2488; // @[LoadQueue.scala 96:50:@5801.6]
  assign _T_2491 = _T_2489 == 1'h0; // @[LoadQueue.scala 96:34:@5802.6]
  assign _T_2493 = previousStoreHead <= offsetQ_9; // @[LoadQueue.scala 101:36:@5810.8]
  assign _T_2494 = offsetQ_9 < io_storeHead; // @[LoadQueue.scala 101:86:@5811.8]
  assign _T_2495 = _T_2493 & _T_2494; // @[LoadQueue.scala 101:61:@5812.8]
  assign _T_2498 = io_storeHead <= offsetQ_9; // @[LoadQueue.scala 103:69:@5818.10]
  assign _T_2499 = offsetQ_9 < previousStoreHead; // @[LoadQueue.scala 104:31:@5819.10]
  assign _T_2500 = _T_2498 & _T_2499; // @[LoadQueue.scala 103:94:@5820.10]
  assign _T_2502 = _T_2500 == 1'h0; // @[LoadQueue.scala 103:54:@5821.10]
  assign _T_2503 = _T_2227 & _T_2502; // @[LoadQueue.scala 103:51:@5822.10]
  assign _GEN_740 = _T_2503 ? 1'h0 : checkBits_9; // @[LoadQueue.scala 104:53:@5823.10]
  assign _GEN_741 = _T_2495 ? 1'h0 : _GEN_740; // @[LoadQueue.scala 101:102:@5813.8]
  assign _GEN_742 = io_storeEmpty ? 1'h0 : _GEN_741; // @[LoadQueue.scala 99:27:@5806.6]
  assign _GEN_743 = initBits_9 ? _T_2491 : _GEN_742; // @[LoadQueue.scala 95:34:@5791.4]
  assign _T_2516 = _GEN_355 + 4'h1; // @[util.scala 10:8:@5834.6]
  assign _GEN_58 = _T_2516 % 5'h10; // @[util.scala 10:14:@5835.6]
  assign _T_2517 = _GEN_58[4:0]; // @[util.scala 10:14:@5835.6]
  assign _T_2518 = _T_2517 == _GEN_2327; // @[LoadQueue.scala 97:56:@5836.6]
  assign _T_2519 = io_storeEmpty & _T_2518; // @[LoadQueue.scala 96:50:@5837.6]
  assign _T_2521 = _T_2519 == 1'h0; // @[LoadQueue.scala 96:34:@5838.6]
  assign _T_2523 = previousStoreHead <= offsetQ_10; // @[LoadQueue.scala 101:36:@5846.8]
  assign _T_2524 = offsetQ_10 < io_storeHead; // @[LoadQueue.scala 101:86:@5847.8]
  assign _T_2525 = _T_2523 & _T_2524; // @[LoadQueue.scala 101:61:@5848.8]
  assign _T_2528 = io_storeHead <= offsetQ_10; // @[LoadQueue.scala 103:69:@5854.10]
  assign _T_2529 = offsetQ_10 < previousStoreHead; // @[LoadQueue.scala 104:31:@5855.10]
  assign _T_2530 = _T_2528 & _T_2529; // @[LoadQueue.scala 103:94:@5856.10]
  assign _T_2532 = _T_2530 == 1'h0; // @[LoadQueue.scala 103:54:@5857.10]
  assign _T_2533 = _T_2227 & _T_2532; // @[LoadQueue.scala 103:51:@5858.10]
  assign _GEN_760 = _T_2533 ? 1'h0 : checkBits_10; // @[LoadQueue.scala 104:53:@5859.10]
  assign _GEN_761 = _T_2525 ? 1'h0 : _GEN_760; // @[LoadQueue.scala 101:102:@5849.8]
  assign _GEN_762 = io_storeEmpty ? 1'h0 : _GEN_761; // @[LoadQueue.scala 99:27:@5842.6]
  assign _GEN_763 = initBits_10 ? _T_2521 : _GEN_762; // @[LoadQueue.scala 95:34:@5827.4]
  assign _T_2546 = _GEN_389 + 4'h1; // @[util.scala 10:8:@5870.6]
  assign _GEN_59 = _T_2546 % 5'h10; // @[util.scala 10:14:@5871.6]
  assign _T_2547 = _GEN_59[4:0]; // @[util.scala 10:14:@5871.6]
  assign _T_2548 = _T_2547 == _GEN_2327; // @[LoadQueue.scala 97:56:@5872.6]
  assign _T_2549 = io_storeEmpty & _T_2548; // @[LoadQueue.scala 96:50:@5873.6]
  assign _T_2551 = _T_2549 == 1'h0; // @[LoadQueue.scala 96:34:@5874.6]
  assign _T_2553 = previousStoreHead <= offsetQ_11; // @[LoadQueue.scala 101:36:@5882.8]
  assign _T_2554 = offsetQ_11 < io_storeHead; // @[LoadQueue.scala 101:86:@5883.8]
  assign _T_2555 = _T_2553 & _T_2554; // @[LoadQueue.scala 101:61:@5884.8]
  assign _T_2558 = io_storeHead <= offsetQ_11; // @[LoadQueue.scala 103:69:@5890.10]
  assign _T_2559 = offsetQ_11 < previousStoreHead; // @[LoadQueue.scala 104:31:@5891.10]
  assign _T_2560 = _T_2558 & _T_2559; // @[LoadQueue.scala 103:94:@5892.10]
  assign _T_2562 = _T_2560 == 1'h0; // @[LoadQueue.scala 103:54:@5893.10]
  assign _T_2563 = _T_2227 & _T_2562; // @[LoadQueue.scala 103:51:@5894.10]
  assign _GEN_780 = _T_2563 ? 1'h0 : checkBits_11; // @[LoadQueue.scala 104:53:@5895.10]
  assign _GEN_781 = _T_2555 ? 1'h0 : _GEN_780; // @[LoadQueue.scala 101:102:@5885.8]
  assign _GEN_782 = io_storeEmpty ? 1'h0 : _GEN_781; // @[LoadQueue.scala 99:27:@5878.6]
  assign _GEN_783 = initBits_11 ? _T_2551 : _GEN_782; // @[LoadQueue.scala 95:34:@5863.4]
  assign _T_2576 = _GEN_423 + 4'h1; // @[util.scala 10:8:@5906.6]
  assign _GEN_60 = _T_2576 % 5'h10; // @[util.scala 10:14:@5907.6]
  assign _T_2577 = _GEN_60[4:0]; // @[util.scala 10:14:@5907.6]
  assign _T_2578 = _T_2577 == _GEN_2327; // @[LoadQueue.scala 97:56:@5908.6]
  assign _T_2579 = io_storeEmpty & _T_2578; // @[LoadQueue.scala 96:50:@5909.6]
  assign _T_2581 = _T_2579 == 1'h0; // @[LoadQueue.scala 96:34:@5910.6]
  assign _T_2583 = previousStoreHead <= offsetQ_12; // @[LoadQueue.scala 101:36:@5918.8]
  assign _T_2584 = offsetQ_12 < io_storeHead; // @[LoadQueue.scala 101:86:@5919.8]
  assign _T_2585 = _T_2583 & _T_2584; // @[LoadQueue.scala 101:61:@5920.8]
  assign _T_2588 = io_storeHead <= offsetQ_12; // @[LoadQueue.scala 103:69:@5926.10]
  assign _T_2589 = offsetQ_12 < previousStoreHead; // @[LoadQueue.scala 104:31:@5927.10]
  assign _T_2590 = _T_2588 & _T_2589; // @[LoadQueue.scala 103:94:@5928.10]
  assign _T_2592 = _T_2590 == 1'h0; // @[LoadQueue.scala 103:54:@5929.10]
  assign _T_2593 = _T_2227 & _T_2592; // @[LoadQueue.scala 103:51:@5930.10]
  assign _GEN_800 = _T_2593 ? 1'h0 : checkBits_12; // @[LoadQueue.scala 104:53:@5931.10]
  assign _GEN_801 = _T_2585 ? 1'h0 : _GEN_800; // @[LoadQueue.scala 101:102:@5921.8]
  assign _GEN_802 = io_storeEmpty ? 1'h0 : _GEN_801; // @[LoadQueue.scala 99:27:@5914.6]
  assign _GEN_803 = initBits_12 ? _T_2581 : _GEN_802; // @[LoadQueue.scala 95:34:@5899.4]
  assign _T_2606 = _GEN_457 + 4'h1; // @[util.scala 10:8:@5942.6]
  assign _GEN_61 = _T_2606 % 5'h10; // @[util.scala 10:14:@5943.6]
  assign _T_2607 = _GEN_61[4:0]; // @[util.scala 10:14:@5943.6]
  assign _T_2608 = _T_2607 == _GEN_2327; // @[LoadQueue.scala 97:56:@5944.6]
  assign _T_2609 = io_storeEmpty & _T_2608; // @[LoadQueue.scala 96:50:@5945.6]
  assign _T_2611 = _T_2609 == 1'h0; // @[LoadQueue.scala 96:34:@5946.6]
  assign _T_2613 = previousStoreHead <= offsetQ_13; // @[LoadQueue.scala 101:36:@5954.8]
  assign _T_2614 = offsetQ_13 < io_storeHead; // @[LoadQueue.scala 101:86:@5955.8]
  assign _T_2615 = _T_2613 & _T_2614; // @[LoadQueue.scala 101:61:@5956.8]
  assign _T_2618 = io_storeHead <= offsetQ_13; // @[LoadQueue.scala 103:69:@5962.10]
  assign _T_2619 = offsetQ_13 < previousStoreHead; // @[LoadQueue.scala 104:31:@5963.10]
  assign _T_2620 = _T_2618 & _T_2619; // @[LoadQueue.scala 103:94:@5964.10]
  assign _T_2622 = _T_2620 == 1'h0; // @[LoadQueue.scala 103:54:@5965.10]
  assign _T_2623 = _T_2227 & _T_2622; // @[LoadQueue.scala 103:51:@5966.10]
  assign _GEN_820 = _T_2623 ? 1'h0 : checkBits_13; // @[LoadQueue.scala 104:53:@5967.10]
  assign _GEN_821 = _T_2615 ? 1'h0 : _GEN_820; // @[LoadQueue.scala 101:102:@5957.8]
  assign _GEN_822 = io_storeEmpty ? 1'h0 : _GEN_821; // @[LoadQueue.scala 99:27:@5950.6]
  assign _GEN_823 = initBits_13 ? _T_2611 : _GEN_822; // @[LoadQueue.scala 95:34:@5935.4]
  assign _T_2636 = _GEN_491 + 4'h1; // @[util.scala 10:8:@5978.6]
  assign _GEN_62 = _T_2636 % 5'h10; // @[util.scala 10:14:@5979.6]
  assign _T_2637 = _GEN_62[4:0]; // @[util.scala 10:14:@5979.6]
  assign _T_2638 = _T_2637 == _GEN_2327; // @[LoadQueue.scala 97:56:@5980.6]
  assign _T_2639 = io_storeEmpty & _T_2638; // @[LoadQueue.scala 96:50:@5981.6]
  assign _T_2641 = _T_2639 == 1'h0; // @[LoadQueue.scala 96:34:@5982.6]
  assign _T_2643 = previousStoreHead <= offsetQ_14; // @[LoadQueue.scala 101:36:@5990.8]
  assign _T_2644 = offsetQ_14 < io_storeHead; // @[LoadQueue.scala 101:86:@5991.8]
  assign _T_2645 = _T_2643 & _T_2644; // @[LoadQueue.scala 101:61:@5992.8]
  assign _T_2648 = io_storeHead <= offsetQ_14; // @[LoadQueue.scala 103:69:@5998.10]
  assign _T_2649 = offsetQ_14 < previousStoreHead; // @[LoadQueue.scala 104:31:@5999.10]
  assign _T_2650 = _T_2648 & _T_2649; // @[LoadQueue.scala 103:94:@6000.10]
  assign _T_2652 = _T_2650 == 1'h0; // @[LoadQueue.scala 103:54:@6001.10]
  assign _T_2653 = _T_2227 & _T_2652; // @[LoadQueue.scala 103:51:@6002.10]
  assign _GEN_840 = _T_2653 ? 1'h0 : checkBits_14; // @[LoadQueue.scala 104:53:@6003.10]
  assign _GEN_841 = _T_2645 ? 1'h0 : _GEN_840; // @[LoadQueue.scala 101:102:@5993.8]
  assign _GEN_842 = io_storeEmpty ? 1'h0 : _GEN_841; // @[LoadQueue.scala 99:27:@5986.6]
  assign _GEN_843 = initBits_14 ? _T_2641 : _GEN_842; // @[LoadQueue.scala 95:34:@5971.4]
  assign _T_2666 = _GEN_525 + 4'h1; // @[util.scala 10:8:@6014.6]
  assign _GEN_63 = _T_2666 % 5'h10; // @[util.scala 10:14:@6015.6]
  assign _T_2667 = _GEN_63[4:0]; // @[util.scala 10:14:@6015.6]
  assign _T_2668 = _T_2667 == _GEN_2327; // @[LoadQueue.scala 97:56:@6016.6]
  assign _T_2669 = io_storeEmpty & _T_2668; // @[LoadQueue.scala 96:50:@6017.6]
  assign _T_2671 = _T_2669 == 1'h0; // @[LoadQueue.scala 96:34:@6018.6]
  assign _T_2673 = previousStoreHead <= offsetQ_15; // @[LoadQueue.scala 101:36:@6026.8]
  assign _T_2674 = offsetQ_15 < io_storeHead; // @[LoadQueue.scala 101:86:@6027.8]
  assign _T_2675 = _T_2673 & _T_2674; // @[LoadQueue.scala 101:61:@6028.8]
  assign _T_2678 = io_storeHead <= offsetQ_15; // @[LoadQueue.scala 103:69:@6034.10]
  assign _T_2679 = offsetQ_15 < previousStoreHead; // @[LoadQueue.scala 104:31:@6035.10]
  assign _T_2680 = _T_2678 & _T_2679; // @[LoadQueue.scala 103:94:@6036.10]
  assign _T_2682 = _T_2680 == 1'h0; // @[LoadQueue.scala 103:54:@6037.10]
  assign _T_2683 = _T_2227 & _T_2682; // @[LoadQueue.scala 103:51:@6038.10]
  assign _GEN_860 = _T_2683 ? 1'h0 : checkBits_15; // @[LoadQueue.scala 104:53:@6039.10]
  assign _GEN_861 = _T_2675 ? 1'h0 : _GEN_860; // @[LoadQueue.scala 101:102:@6029.8]
  assign _GEN_862 = io_storeEmpty ? 1'h0 : _GEN_861; // @[LoadQueue.scala 99:27:@6022.6]
  assign _GEN_863 = initBits_15 ? _T_2671 : _GEN_862; // @[LoadQueue.scala 95:34:@6007.4]
  assign _T_2687 = 16'h1 << io_storeHead; // @[OneHot.scala 52:12:@6044.4]
  assign _T_2689 = _T_2687[0]; // @[util.scala 60:60:@6046.4]
  assign _T_2690 = _T_2687[1]; // @[util.scala 60:60:@6047.4]
  assign _T_2691 = _T_2687[2]; // @[util.scala 60:60:@6048.4]
  assign _T_2692 = _T_2687[3]; // @[util.scala 60:60:@6049.4]
  assign _T_2693 = _T_2687[4]; // @[util.scala 60:60:@6050.4]
  assign _T_2694 = _T_2687[5]; // @[util.scala 60:60:@6051.4]
  assign _T_2695 = _T_2687[6]; // @[util.scala 60:60:@6052.4]
  assign _T_2696 = _T_2687[7]; // @[util.scala 60:60:@6053.4]
  assign _T_2697 = _T_2687[8]; // @[util.scala 60:60:@6054.4]
  assign _T_2698 = _T_2687[9]; // @[util.scala 60:60:@6055.4]
  assign _T_2699 = _T_2687[10]; // @[util.scala 60:60:@6056.4]
  assign _T_2700 = _T_2687[11]; // @[util.scala 60:60:@6057.4]
  assign _T_2701 = _T_2687[12]; // @[util.scala 60:60:@6058.4]
  assign _T_2702 = _T_2687[13]; // @[util.scala 60:60:@6059.4]
  assign _T_2703 = _T_2687[14]; // @[util.scala 60:60:@6060.4]
  assign _T_2704 = _T_2687[15]; // @[util.scala 60:60:@6061.4]
  assign _T_4835 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@7585.4]
  assign _T_4842 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8}; // @[Mux.scala 19:72:@7592.4]
  assign _T_4843 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,_T_4835}; // @[Mux.scala 19:72:@7593.4]
  assign _T_4845 = _T_2689 ? _T_4843 : 512'h0; // @[Mux.scala 19:72:@7594.4]
  assign _T_4852 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@7601.4]
  assign _T_4859 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9}; // @[Mux.scala 19:72:@7608.4]
  assign _T_4860 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,_T_4852}; // @[Mux.scala 19:72:@7609.4]
  assign _T_4862 = _T_2690 ? _T_4860 : 512'h0; // @[Mux.scala 19:72:@7610.4]
  assign _T_4869 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@7617.4]
  assign _T_4876 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10}; // @[Mux.scala 19:72:@7624.4]
  assign _T_4877 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,_T_4869}; // @[Mux.scala 19:72:@7625.4]
  assign _T_4879 = _T_2691 ? _T_4877 : 512'h0; // @[Mux.scala 19:72:@7626.4]
  assign _T_4886 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@7633.4]
  assign _T_4893 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11}; // @[Mux.scala 19:72:@7640.4]
  assign _T_4894 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,_T_4886}; // @[Mux.scala 19:72:@7641.4]
  assign _T_4896 = _T_2692 ? _T_4894 : 512'h0; // @[Mux.scala 19:72:@7642.4]
  assign _T_4903 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@7649.4]
  assign _T_4910 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12}; // @[Mux.scala 19:72:@7656.4]
  assign _T_4911 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,_T_4903}; // @[Mux.scala 19:72:@7657.4]
  assign _T_4913 = _T_2693 ? _T_4911 : 512'h0; // @[Mux.scala 19:72:@7658.4]
  assign _T_4920 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@7665.4]
  assign _T_4927 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13}; // @[Mux.scala 19:72:@7672.4]
  assign _T_4928 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,_T_4920}; // @[Mux.scala 19:72:@7673.4]
  assign _T_4930 = _T_2694 ? _T_4928 : 512'h0; // @[Mux.scala 19:72:@7674.4]
  assign _T_4937 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@7681.4]
  assign _T_4944 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14}; // @[Mux.scala 19:72:@7688.4]
  assign _T_4945 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,_T_4937}; // @[Mux.scala 19:72:@7689.4]
  assign _T_4947 = _T_2695 ? _T_4945 : 512'h0; // @[Mux.scala 19:72:@7690.4]
  assign _T_4954 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7}; // @[Mux.scala 19:72:@7697.4]
  assign _T_4961 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15}; // @[Mux.scala 19:72:@7704.4]
  assign _T_4962 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,_T_4954}; // @[Mux.scala 19:72:@7705.4]
  assign _T_4964 = _T_2696 ? _T_4962 : 512'h0; // @[Mux.scala 19:72:@7706.4]
  assign _T_4979 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,_T_4842}; // @[Mux.scala 19:72:@7721.4]
  assign _T_4981 = _T_2697 ? _T_4979 : 512'h0; // @[Mux.scala 19:72:@7722.4]
  assign _T_4996 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,_T_4859}; // @[Mux.scala 19:72:@7737.4]
  assign _T_4998 = _T_2698 ? _T_4996 : 512'h0; // @[Mux.scala 19:72:@7738.4]
  assign _T_5013 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,_T_4876}; // @[Mux.scala 19:72:@7753.4]
  assign _T_5015 = _T_2699 ? _T_5013 : 512'h0; // @[Mux.scala 19:72:@7754.4]
  assign _T_5030 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,_T_4893}; // @[Mux.scala 19:72:@7769.4]
  assign _T_5032 = _T_2700 ? _T_5030 : 512'h0; // @[Mux.scala 19:72:@7770.4]
  assign _T_5047 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,_T_4910}; // @[Mux.scala 19:72:@7785.4]
  assign _T_5049 = _T_2701 ? _T_5047 : 512'h0; // @[Mux.scala 19:72:@7786.4]
  assign _T_5064 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,_T_4927}; // @[Mux.scala 19:72:@7801.4]
  assign _T_5066 = _T_2702 ? _T_5064 : 512'h0; // @[Mux.scala 19:72:@7802.4]
  assign _T_5081 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,_T_4944}; // @[Mux.scala 19:72:@7817.4]
  assign _T_5083 = _T_2703 ? _T_5081 : 512'h0; // @[Mux.scala 19:72:@7818.4]
  assign _T_5098 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,_T_4961}; // @[Mux.scala 19:72:@7833.4]
  assign _T_5100 = _T_2704 ? _T_5098 : 512'h0; // @[Mux.scala 19:72:@7834.4]
  assign _T_5101 = _T_4845 | _T_4862; // @[Mux.scala 19:72:@7835.4]
  assign _T_5102 = _T_5101 | _T_4879; // @[Mux.scala 19:72:@7836.4]
  assign _T_5103 = _T_5102 | _T_4896; // @[Mux.scala 19:72:@7837.4]
  assign _T_5104 = _T_5103 | _T_4913; // @[Mux.scala 19:72:@7838.4]
  assign _T_5105 = _T_5104 | _T_4930; // @[Mux.scala 19:72:@7839.4]
  assign _T_5106 = _T_5105 | _T_4947; // @[Mux.scala 19:72:@7840.4]
  assign _T_5107 = _T_5106 | _T_4964; // @[Mux.scala 19:72:@7841.4]
  assign _T_5108 = _T_5107 | _T_4981; // @[Mux.scala 19:72:@7842.4]
  assign _T_5109 = _T_5108 | _T_4998; // @[Mux.scala 19:72:@7843.4]
  assign _T_5110 = _T_5109 | _T_5015; // @[Mux.scala 19:72:@7844.4]
  assign _T_5111 = _T_5110 | _T_5032; // @[Mux.scala 19:72:@7845.4]
  assign _T_5112 = _T_5111 | _T_5049; // @[Mux.scala 19:72:@7846.4]
  assign _T_5113 = _T_5112 | _T_5066; // @[Mux.scala 19:72:@7847.4]
  assign _T_5114 = _T_5113 | _T_5083; // @[Mux.scala 19:72:@7848.4]
  assign _T_5115 = _T_5114 | _T_5100; // @[Mux.scala 19:72:@7849.4]
  assign _T_5692 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@8199.4]
  assign _T_5699 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8}; // @[Mux.scala 19:72:@8206.4]
  assign _T_5700 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,_T_5692}; // @[Mux.scala 19:72:@8207.4]
  assign _T_5702 = _T_2689 ? _T_5700 : 16'h0; // @[Mux.scala 19:72:@8208.4]
  assign _T_5709 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@8215.4]
  assign _T_5716 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9}; // @[Mux.scala 19:72:@8222.4]
  assign _T_5717 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,_T_5709}; // @[Mux.scala 19:72:@8223.4]
  assign _T_5719 = _T_2690 ? _T_5717 : 16'h0; // @[Mux.scala 19:72:@8224.4]
  assign _T_5726 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@8231.4]
  assign _T_5733 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10}; // @[Mux.scala 19:72:@8238.4]
  assign _T_5734 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,_T_5726}; // @[Mux.scala 19:72:@8239.4]
  assign _T_5736 = _T_2691 ? _T_5734 : 16'h0; // @[Mux.scala 19:72:@8240.4]
  assign _T_5743 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@8247.4]
  assign _T_5750 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11}; // @[Mux.scala 19:72:@8254.4]
  assign _T_5751 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,_T_5743}; // @[Mux.scala 19:72:@8255.4]
  assign _T_5753 = _T_2692 ? _T_5751 : 16'h0; // @[Mux.scala 19:72:@8256.4]
  assign _T_5760 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@8263.4]
  assign _T_5767 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12}; // @[Mux.scala 19:72:@8270.4]
  assign _T_5768 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,_T_5760}; // @[Mux.scala 19:72:@8271.4]
  assign _T_5770 = _T_2693 ? _T_5768 : 16'h0; // @[Mux.scala 19:72:@8272.4]
  assign _T_5777 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@8279.4]
  assign _T_5784 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13}; // @[Mux.scala 19:72:@8286.4]
  assign _T_5785 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,_T_5777}; // @[Mux.scala 19:72:@8287.4]
  assign _T_5787 = _T_2694 ? _T_5785 : 16'h0; // @[Mux.scala 19:72:@8288.4]
  assign _T_5794 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@8295.4]
  assign _T_5801 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14}; // @[Mux.scala 19:72:@8302.4]
  assign _T_5802 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,_T_5794}; // @[Mux.scala 19:72:@8303.4]
  assign _T_5804 = _T_2695 ? _T_5802 : 16'h0; // @[Mux.scala 19:72:@8304.4]
  assign _T_5811 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7}; // @[Mux.scala 19:72:@8311.4]
  assign _T_5818 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15}; // @[Mux.scala 19:72:@8318.4]
  assign _T_5819 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,_T_5811}; // @[Mux.scala 19:72:@8319.4]
  assign _T_5821 = _T_2696 ? _T_5819 : 16'h0; // @[Mux.scala 19:72:@8320.4]
  assign _T_5836 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,_T_5699}; // @[Mux.scala 19:72:@8335.4]
  assign _T_5838 = _T_2697 ? _T_5836 : 16'h0; // @[Mux.scala 19:72:@8336.4]
  assign _T_5853 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,_T_5716}; // @[Mux.scala 19:72:@8351.4]
  assign _T_5855 = _T_2698 ? _T_5853 : 16'h0; // @[Mux.scala 19:72:@8352.4]
  assign _T_5870 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,_T_5733}; // @[Mux.scala 19:72:@8367.4]
  assign _T_5872 = _T_2699 ? _T_5870 : 16'h0; // @[Mux.scala 19:72:@8368.4]
  assign _T_5887 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,_T_5750}; // @[Mux.scala 19:72:@8383.4]
  assign _T_5889 = _T_2700 ? _T_5887 : 16'h0; // @[Mux.scala 19:72:@8384.4]
  assign _T_5904 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,_T_5767}; // @[Mux.scala 19:72:@8399.4]
  assign _T_5906 = _T_2701 ? _T_5904 : 16'h0; // @[Mux.scala 19:72:@8400.4]
  assign _T_5921 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,_T_5784}; // @[Mux.scala 19:72:@8415.4]
  assign _T_5923 = _T_2702 ? _T_5921 : 16'h0; // @[Mux.scala 19:72:@8416.4]
  assign _T_5938 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,_T_5801}; // @[Mux.scala 19:72:@8431.4]
  assign _T_5940 = _T_2703 ? _T_5938 : 16'h0; // @[Mux.scala 19:72:@8432.4]
  assign _T_5955 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,_T_5818}; // @[Mux.scala 19:72:@8447.4]
  assign _T_5957 = _T_2704 ? _T_5955 : 16'h0; // @[Mux.scala 19:72:@8448.4]
  assign _T_5958 = _T_5702 | _T_5719; // @[Mux.scala 19:72:@8449.4]
  assign _T_5959 = _T_5958 | _T_5736; // @[Mux.scala 19:72:@8450.4]
  assign _T_5960 = _T_5959 | _T_5753; // @[Mux.scala 19:72:@8451.4]
  assign _T_5961 = _T_5960 | _T_5770; // @[Mux.scala 19:72:@8452.4]
  assign _T_5962 = _T_5961 | _T_5787; // @[Mux.scala 19:72:@8453.4]
  assign _T_5963 = _T_5962 | _T_5804; // @[Mux.scala 19:72:@8454.4]
  assign _T_5964 = _T_5963 | _T_5821; // @[Mux.scala 19:72:@8455.4]
  assign _T_5965 = _T_5964 | _T_5838; // @[Mux.scala 19:72:@8456.4]
  assign _T_5966 = _T_5965 | _T_5855; // @[Mux.scala 19:72:@8457.4]
  assign _T_5967 = _T_5966 | _T_5872; // @[Mux.scala 19:72:@8458.4]
  assign _T_5968 = _T_5967 | _T_5889; // @[Mux.scala 19:72:@8459.4]
  assign _T_5969 = _T_5968 | _T_5906; // @[Mux.scala 19:72:@8460.4]
  assign _T_5970 = _T_5969 | _T_5923; // @[Mux.scala 19:72:@8461.4]
  assign _T_5971 = _T_5970 | _T_5940; // @[Mux.scala 19:72:@8462.4]
  assign _T_5972 = _T_5971 | _T_5957; // @[Mux.scala 19:72:@8463.4]
  assign _T_6113 = io_storeHead < io_storeTail; // @[LoadQueue.scala 121:105:@8499.4]
  assign _T_6115 = io_storeHead <= 4'h0; // @[LoadQueue.scala 122:18:@8500.4]
  assign _T_6117 = 4'h0 < io_storeTail; // @[LoadQueue.scala 122:36:@8501.4]
  assign _T_6118 = _T_6115 & _T_6117; // @[LoadQueue.scala 122:27:@8502.4]
  assign _T_6120 = io_storeEmpty == 1'h0; // @[LoadQueue.scala 122:52:@8503.4]
  assign _T_6122 = io_storeTail <= 4'h0; // @[LoadQueue.scala 122:85:@8504.4]
  assign _T_6124 = 4'h0 < io_storeHead; // @[LoadQueue.scala 122:103:@8505.4]
  assign _T_6125 = _T_6122 & _T_6124; // @[LoadQueue.scala 122:94:@8506.4]
  assign _T_6127 = _T_6125 == 1'h0; // @[LoadQueue.scala 122:70:@8507.4]
  assign _T_6128 = _T_6120 & _T_6127; // @[LoadQueue.scala 122:67:@8508.4]
  assign validEntriesInStoreQ_0 = _T_6113 ? _T_6118 : _T_6128; // @[LoadQueue.scala 121:91:@8509.4]
  assign _T_6132 = io_storeHead <= 4'h1; // @[LoadQueue.scala 122:18:@8511.4]
  assign _T_6134 = 4'h1 < io_storeTail; // @[LoadQueue.scala 122:36:@8512.4]
  assign _T_6135 = _T_6132 & _T_6134; // @[LoadQueue.scala 122:27:@8513.4]
  assign _T_6139 = io_storeTail <= 4'h1; // @[LoadQueue.scala 122:85:@8515.4]
  assign _T_6141 = 4'h1 < io_storeHead; // @[LoadQueue.scala 122:103:@8516.4]
  assign _T_6142 = _T_6139 & _T_6141; // @[LoadQueue.scala 122:94:@8517.4]
  assign _T_6144 = _T_6142 == 1'h0; // @[LoadQueue.scala 122:70:@8518.4]
  assign _T_6145 = _T_6120 & _T_6144; // @[LoadQueue.scala 122:67:@8519.4]
  assign validEntriesInStoreQ_1 = _T_6113 ? _T_6135 : _T_6145; // @[LoadQueue.scala 121:91:@8520.4]
  assign _T_6149 = io_storeHead <= 4'h2; // @[LoadQueue.scala 122:18:@8522.4]
  assign _T_6151 = 4'h2 < io_storeTail; // @[LoadQueue.scala 122:36:@8523.4]
  assign _T_6152 = _T_6149 & _T_6151; // @[LoadQueue.scala 122:27:@8524.4]
  assign _T_6156 = io_storeTail <= 4'h2; // @[LoadQueue.scala 122:85:@8526.4]
  assign _T_6158 = 4'h2 < io_storeHead; // @[LoadQueue.scala 122:103:@8527.4]
  assign _T_6159 = _T_6156 & _T_6158; // @[LoadQueue.scala 122:94:@8528.4]
  assign _T_6161 = _T_6159 == 1'h0; // @[LoadQueue.scala 122:70:@8529.4]
  assign _T_6162 = _T_6120 & _T_6161; // @[LoadQueue.scala 122:67:@8530.4]
  assign validEntriesInStoreQ_2 = _T_6113 ? _T_6152 : _T_6162; // @[LoadQueue.scala 121:91:@8531.4]
  assign _T_6166 = io_storeHead <= 4'h3; // @[LoadQueue.scala 122:18:@8533.4]
  assign _T_6168 = 4'h3 < io_storeTail; // @[LoadQueue.scala 122:36:@8534.4]
  assign _T_6169 = _T_6166 & _T_6168; // @[LoadQueue.scala 122:27:@8535.4]
  assign _T_6173 = io_storeTail <= 4'h3; // @[LoadQueue.scala 122:85:@8537.4]
  assign _T_6175 = 4'h3 < io_storeHead; // @[LoadQueue.scala 122:103:@8538.4]
  assign _T_6176 = _T_6173 & _T_6175; // @[LoadQueue.scala 122:94:@8539.4]
  assign _T_6178 = _T_6176 == 1'h0; // @[LoadQueue.scala 122:70:@8540.4]
  assign _T_6179 = _T_6120 & _T_6178; // @[LoadQueue.scala 122:67:@8541.4]
  assign validEntriesInStoreQ_3 = _T_6113 ? _T_6169 : _T_6179; // @[LoadQueue.scala 121:91:@8542.4]
  assign _T_6183 = io_storeHead <= 4'h4; // @[LoadQueue.scala 122:18:@8544.4]
  assign _T_6185 = 4'h4 < io_storeTail; // @[LoadQueue.scala 122:36:@8545.4]
  assign _T_6186 = _T_6183 & _T_6185; // @[LoadQueue.scala 122:27:@8546.4]
  assign _T_6190 = io_storeTail <= 4'h4; // @[LoadQueue.scala 122:85:@8548.4]
  assign _T_6192 = 4'h4 < io_storeHead; // @[LoadQueue.scala 122:103:@8549.4]
  assign _T_6193 = _T_6190 & _T_6192; // @[LoadQueue.scala 122:94:@8550.4]
  assign _T_6195 = _T_6193 == 1'h0; // @[LoadQueue.scala 122:70:@8551.4]
  assign _T_6196 = _T_6120 & _T_6195; // @[LoadQueue.scala 122:67:@8552.4]
  assign validEntriesInStoreQ_4 = _T_6113 ? _T_6186 : _T_6196; // @[LoadQueue.scala 121:91:@8553.4]
  assign _T_6200 = io_storeHead <= 4'h5; // @[LoadQueue.scala 122:18:@8555.4]
  assign _T_6202 = 4'h5 < io_storeTail; // @[LoadQueue.scala 122:36:@8556.4]
  assign _T_6203 = _T_6200 & _T_6202; // @[LoadQueue.scala 122:27:@8557.4]
  assign _T_6207 = io_storeTail <= 4'h5; // @[LoadQueue.scala 122:85:@8559.4]
  assign _T_6209 = 4'h5 < io_storeHead; // @[LoadQueue.scala 122:103:@8560.4]
  assign _T_6210 = _T_6207 & _T_6209; // @[LoadQueue.scala 122:94:@8561.4]
  assign _T_6212 = _T_6210 == 1'h0; // @[LoadQueue.scala 122:70:@8562.4]
  assign _T_6213 = _T_6120 & _T_6212; // @[LoadQueue.scala 122:67:@8563.4]
  assign validEntriesInStoreQ_5 = _T_6113 ? _T_6203 : _T_6213; // @[LoadQueue.scala 121:91:@8564.4]
  assign _T_6217 = io_storeHead <= 4'h6; // @[LoadQueue.scala 122:18:@8566.4]
  assign _T_6219 = 4'h6 < io_storeTail; // @[LoadQueue.scala 122:36:@8567.4]
  assign _T_6220 = _T_6217 & _T_6219; // @[LoadQueue.scala 122:27:@8568.4]
  assign _T_6224 = io_storeTail <= 4'h6; // @[LoadQueue.scala 122:85:@8570.4]
  assign _T_6226 = 4'h6 < io_storeHead; // @[LoadQueue.scala 122:103:@8571.4]
  assign _T_6227 = _T_6224 & _T_6226; // @[LoadQueue.scala 122:94:@8572.4]
  assign _T_6229 = _T_6227 == 1'h0; // @[LoadQueue.scala 122:70:@8573.4]
  assign _T_6230 = _T_6120 & _T_6229; // @[LoadQueue.scala 122:67:@8574.4]
  assign validEntriesInStoreQ_6 = _T_6113 ? _T_6220 : _T_6230; // @[LoadQueue.scala 121:91:@8575.4]
  assign _T_6234 = io_storeHead <= 4'h7; // @[LoadQueue.scala 122:18:@8577.4]
  assign _T_6236 = 4'h7 < io_storeTail; // @[LoadQueue.scala 122:36:@8578.4]
  assign _T_6237 = _T_6234 & _T_6236; // @[LoadQueue.scala 122:27:@8579.4]
  assign _T_6241 = io_storeTail <= 4'h7; // @[LoadQueue.scala 122:85:@8581.4]
  assign _T_6243 = 4'h7 < io_storeHead; // @[LoadQueue.scala 122:103:@8582.4]
  assign _T_6244 = _T_6241 & _T_6243; // @[LoadQueue.scala 122:94:@8583.4]
  assign _T_6246 = _T_6244 == 1'h0; // @[LoadQueue.scala 122:70:@8584.4]
  assign _T_6247 = _T_6120 & _T_6246; // @[LoadQueue.scala 122:67:@8585.4]
  assign validEntriesInStoreQ_7 = _T_6113 ? _T_6237 : _T_6247; // @[LoadQueue.scala 121:91:@8586.4]
  assign _T_6251 = io_storeHead <= 4'h8; // @[LoadQueue.scala 122:18:@8588.4]
  assign _T_6253 = 4'h8 < io_storeTail; // @[LoadQueue.scala 122:36:@8589.4]
  assign _T_6254 = _T_6251 & _T_6253; // @[LoadQueue.scala 122:27:@8590.4]
  assign _T_6258 = io_storeTail <= 4'h8; // @[LoadQueue.scala 122:85:@8592.4]
  assign _T_6260 = 4'h8 < io_storeHead; // @[LoadQueue.scala 122:103:@8593.4]
  assign _T_6261 = _T_6258 & _T_6260; // @[LoadQueue.scala 122:94:@8594.4]
  assign _T_6263 = _T_6261 == 1'h0; // @[LoadQueue.scala 122:70:@8595.4]
  assign _T_6264 = _T_6120 & _T_6263; // @[LoadQueue.scala 122:67:@8596.4]
  assign validEntriesInStoreQ_8 = _T_6113 ? _T_6254 : _T_6264; // @[LoadQueue.scala 121:91:@8597.4]
  assign _T_6268 = io_storeHead <= 4'h9; // @[LoadQueue.scala 122:18:@8599.4]
  assign _T_6270 = 4'h9 < io_storeTail; // @[LoadQueue.scala 122:36:@8600.4]
  assign _T_6271 = _T_6268 & _T_6270; // @[LoadQueue.scala 122:27:@8601.4]
  assign _T_6275 = io_storeTail <= 4'h9; // @[LoadQueue.scala 122:85:@8603.4]
  assign _T_6277 = 4'h9 < io_storeHead; // @[LoadQueue.scala 122:103:@8604.4]
  assign _T_6278 = _T_6275 & _T_6277; // @[LoadQueue.scala 122:94:@8605.4]
  assign _T_6280 = _T_6278 == 1'h0; // @[LoadQueue.scala 122:70:@8606.4]
  assign _T_6281 = _T_6120 & _T_6280; // @[LoadQueue.scala 122:67:@8607.4]
  assign validEntriesInStoreQ_9 = _T_6113 ? _T_6271 : _T_6281; // @[LoadQueue.scala 121:91:@8608.4]
  assign _T_6285 = io_storeHead <= 4'ha; // @[LoadQueue.scala 122:18:@8610.4]
  assign _T_6287 = 4'ha < io_storeTail; // @[LoadQueue.scala 122:36:@8611.4]
  assign _T_6288 = _T_6285 & _T_6287; // @[LoadQueue.scala 122:27:@8612.4]
  assign _T_6292 = io_storeTail <= 4'ha; // @[LoadQueue.scala 122:85:@8614.4]
  assign _T_6294 = 4'ha < io_storeHead; // @[LoadQueue.scala 122:103:@8615.4]
  assign _T_6295 = _T_6292 & _T_6294; // @[LoadQueue.scala 122:94:@8616.4]
  assign _T_6297 = _T_6295 == 1'h0; // @[LoadQueue.scala 122:70:@8617.4]
  assign _T_6298 = _T_6120 & _T_6297; // @[LoadQueue.scala 122:67:@8618.4]
  assign validEntriesInStoreQ_10 = _T_6113 ? _T_6288 : _T_6298; // @[LoadQueue.scala 121:91:@8619.4]
  assign _T_6302 = io_storeHead <= 4'hb; // @[LoadQueue.scala 122:18:@8621.4]
  assign _T_6304 = 4'hb < io_storeTail; // @[LoadQueue.scala 122:36:@8622.4]
  assign _T_6305 = _T_6302 & _T_6304; // @[LoadQueue.scala 122:27:@8623.4]
  assign _T_6309 = io_storeTail <= 4'hb; // @[LoadQueue.scala 122:85:@8625.4]
  assign _T_6311 = 4'hb < io_storeHead; // @[LoadQueue.scala 122:103:@8626.4]
  assign _T_6312 = _T_6309 & _T_6311; // @[LoadQueue.scala 122:94:@8627.4]
  assign _T_6314 = _T_6312 == 1'h0; // @[LoadQueue.scala 122:70:@8628.4]
  assign _T_6315 = _T_6120 & _T_6314; // @[LoadQueue.scala 122:67:@8629.4]
  assign validEntriesInStoreQ_11 = _T_6113 ? _T_6305 : _T_6315; // @[LoadQueue.scala 121:91:@8630.4]
  assign _T_6319 = io_storeHead <= 4'hc; // @[LoadQueue.scala 122:18:@8632.4]
  assign _T_6321 = 4'hc < io_storeTail; // @[LoadQueue.scala 122:36:@8633.4]
  assign _T_6322 = _T_6319 & _T_6321; // @[LoadQueue.scala 122:27:@8634.4]
  assign _T_6326 = io_storeTail <= 4'hc; // @[LoadQueue.scala 122:85:@8636.4]
  assign _T_6328 = 4'hc < io_storeHead; // @[LoadQueue.scala 122:103:@8637.4]
  assign _T_6329 = _T_6326 & _T_6328; // @[LoadQueue.scala 122:94:@8638.4]
  assign _T_6331 = _T_6329 == 1'h0; // @[LoadQueue.scala 122:70:@8639.4]
  assign _T_6332 = _T_6120 & _T_6331; // @[LoadQueue.scala 122:67:@8640.4]
  assign validEntriesInStoreQ_12 = _T_6113 ? _T_6322 : _T_6332; // @[LoadQueue.scala 121:91:@8641.4]
  assign _T_6336 = io_storeHead <= 4'hd; // @[LoadQueue.scala 122:18:@8643.4]
  assign _T_6338 = 4'hd < io_storeTail; // @[LoadQueue.scala 122:36:@8644.4]
  assign _T_6339 = _T_6336 & _T_6338; // @[LoadQueue.scala 122:27:@8645.4]
  assign _T_6343 = io_storeTail <= 4'hd; // @[LoadQueue.scala 122:85:@8647.4]
  assign _T_6345 = 4'hd < io_storeHead; // @[LoadQueue.scala 122:103:@8648.4]
  assign _T_6346 = _T_6343 & _T_6345; // @[LoadQueue.scala 122:94:@8649.4]
  assign _T_6348 = _T_6346 == 1'h0; // @[LoadQueue.scala 122:70:@8650.4]
  assign _T_6349 = _T_6120 & _T_6348; // @[LoadQueue.scala 122:67:@8651.4]
  assign validEntriesInStoreQ_13 = _T_6113 ? _T_6339 : _T_6349; // @[LoadQueue.scala 121:91:@8652.4]
  assign _T_6353 = io_storeHead <= 4'he; // @[LoadQueue.scala 122:18:@8654.4]
  assign _T_6355 = 4'he < io_storeTail; // @[LoadQueue.scala 122:36:@8655.4]
  assign _T_6356 = _T_6353 & _T_6355; // @[LoadQueue.scala 122:27:@8656.4]
  assign _T_6360 = io_storeTail <= 4'he; // @[LoadQueue.scala 122:85:@8658.4]
  assign _T_6362 = 4'he < io_storeHead; // @[LoadQueue.scala 122:103:@8659.4]
  assign _T_6363 = _T_6360 & _T_6362; // @[LoadQueue.scala 122:94:@8660.4]
  assign _T_6365 = _T_6363 == 1'h0; // @[LoadQueue.scala 122:70:@8661.4]
  assign _T_6366 = _T_6120 & _T_6365; // @[LoadQueue.scala 122:67:@8662.4]
  assign validEntriesInStoreQ_14 = _T_6113 ? _T_6356 : _T_6366; // @[LoadQueue.scala 121:91:@8663.4]
  assign validEntriesInStoreQ_15 = _T_6113 ? 1'h0 : _T_6120; // @[LoadQueue.scala 121:91:@8674.4]
  assign storesToCheck_0_0 = _T_2228 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@8701.4]
  assign _T_7654 = 4'h1 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8704.4]
  assign _T_7655 = _T_6132 & _T_7654; // @[LoadQueue.scala 131:72:@8705.4]
  assign _T_7657 = offsetQ_0 < 4'h1; // @[LoadQueue.scala 132:33:@8706.4]
  assign _T_7660 = _T_7657 & _T_6141; // @[LoadQueue.scala 132:41:@8708.4]
  assign _T_7662 = _T_7660 == 1'h0; // @[LoadQueue.scala 132:9:@8709.4]
  assign storesToCheck_0_1 = _T_2228 ? _T_7655 : _T_7662; // @[LoadQueue.scala 131:10:@8710.4]
  assign _T_7668 = 4'h2 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8713.4]
  assign _T_7669 = _T_6149 & _T_7668; // @[LoadQueue.scala 131:72:@8714.4]
  assign _T_7671 = offsetQ_0 < 4'h2; // @[LoadQueue.scala 132:33:@8715.4]
  assign _T_7674 = _T_7671 & _T_6158; // @[LoadQueue.scala 132:41:@8717.4]
  assign _T_7676 = _T_7674 == 1'h0; // @[LoadQueue.scala 132:9:@8718.4]
  assign storesToCheck_0_2 = _T_2228 ? _T_7669 : _T_7676; // @[LoadQueue.scala 131:10:@8719.4]
  assign _T_7682 = 4'h3 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8722.4]
  assign _T_7683 = _T_6166 & _T_7682; // @[LoadQueue.scala 131:72:@8723.4]
  assign _T_7685 = offsetQ_0 < 4'h3; // @[LoadQueue.scala 132:33:@8724.4]
  assign _T_7688 = _T_7685 & _T_6175; // @[LoadQueue.scala 132:41:@8726.4]
  assign _T_7690 = _T_7688 == 1'h0; // @[LoadQueue.scala 132:9:@8727.4]
  assign storesToCheck_0_3 = _T_2228 ? _T_7683 : _T_7690; // @[LoadQueue.scala 131:10:@8728.4]
  assign _T_7696 = 4'h4 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8731.4]
  assign _T_7697 = _T_6183 & _T_7696; // @[LoadQueue.scala 131:72:@8732.4]
  assign _T_7699 = offsetQ_0 < 4'h4; // @[LoadQueue.scala 132:33:@8733.4]
  assign _T_7702 = _T_7699 & _T_6192; // @[LoadQueue.scala 132:41:@8735.4]
  assign _T_7704 = _T_7702 == 1'h0; // @[LoadQueue.scala 132:9:@8736.4]
  assign storesToCheck_0_4 = _T_2228 ? _T_7697 : _T_7704; // @[LoadQueue.scala 131:10:@8737.4]
  assign _T_7710 = 4'h5 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8740.4]
  assign _T_7711 = _T_6200 & _T_7710; // @[LoadQueue.scala 131:72:@8741.4]
  assign _T_7713 = offsetQ_0 < 4'h5; // @[LoadQueue.scala 132:33:@8742.4]
  assign _T_7716 = _T_7713 & _T_6209; // @[LoadQueue.scala 132:41:@8744.4]
  assign _T_7718 = _T_7716 == 1'h0; // @[LoadQueue.scala 132:9:@8745.4]
  assign storesToCheck_0_5 = _T_2228 ? _T_7711 : _T_7718; // @[LoadQueue.scala 131:10:@8746.4]
  assign _T_7724 = 4'h6 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8749.4]
  assign _T_7725 = _T_6217 & _T_7724; // @[LoadQueue.scala 131:72:@8750.4]
  assign _T_7727 = offsetQ_0 < 4'h6; // @[LoadQueue.scala 132:33:@8751.4]
  assign _T_7730 = _T_7727 & _T_6226; // @[LoadQueue.scala 132:41:@8753.4]
  assign _T_7732 = _T_7730 == 1'h0; // @[LoadQueue.scala 132:9:@8754.4]
  assign storesToCheck_0_6 = _T_2228 ? _T_7725 : _T_7732; // @[LoadQueue.scala 131:10:@8755.4]
  assign _T_7738 = 4'h7 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8758.4]
  assign _T_7739 = _T_6234 & _T_7738; // @[LoadQueue.scala 131:72:@8759.4]
  assign _T_7741 = offsetQ_0 < 4'h7; // @[LoadQueue.scala 132:33:@8760.4]
  assign _T_7744 = _T_7741 & _T_6243; // @[LoadQueue.scala 132:41:@8762.4]
  assign _T_7746 = _T_7744 == 1'h0; // @[LoadQueue.scala 132:9:@8763.4]
  assign storesToCheck_0_7 = _T_2228 ? _T_7739 : _T_7746; // @[LoadQueue.scala 131:10:@8764.4]
  assign _T_7752 = 4'h8 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8767.4]
  assign _T_7753 = _T_6251 & _T_7752; // @[LoadQueue.scala 131:72:@8768.4]
  assign _T_7755 = offsetQ_0 < 4'h8; // @[LoadQueue.scala 132:33:@8769.4]
  assign _T_7758 = _T_7755 & _T_6260; // @[LoadQueue.scala 132:41:@8771.4]
  assign _T_7760 = _T_7758 == 1'h0; // @[LoadQueue.scala 132:9:@8772.4]
  assign storesToCheck_0_8 = _T_2228 ? _T_7753 : _T_7760; // @[LoadQueue.scala 131:10:@8773.4]
  assign _T_7766 = 4'h9 <= offsetQ_0; // @[LoadQueue.scala 131:81:@8776.4]
  assign _T_7767 = _T_6268 & _T_7766; // @[LoadQueue.scala 131:72:@8777.4]
  assign _T_7769 = offsetQ_0 < 4'h9; // @[LoadQueue.scala 132:33:@8778.4]
  assign _T_7772 = _T_7769 & _T_6277; // @[LoadQueue.scala 132:41:@8780.4]
  assign _T_7774 = _T_7772 == 1'h0; // @[LoadQueue.scala 132:9:@8781.4]
  assign storesToCheck_0_9 = _T_2228 ? _T_7767 : _T_7774; // @[LoadQueue.scala 131:10:@8782.4]
  assign _T_7780 = 4'ha <= offsetQ_0; // @[LoadQueue.scala 131:81:@8785.4]
  assign _T_7781 = _T_6285 & _T_7780; // @[LoadQueue.scala 131:72:@8786.4]
  assign _T_7783 = offsetQ_0 < 4'ha; // @[LoadQueue.scala 132:33:@8787.4]
  assign _T_7786 = _T_7783 & _T_6294; // @[LoadQueue.scala 132:41:@8789.4]
  assign _T_7788 = _T_7786 == 1'h0; // @[LoadQueue.scala 132:9:@8790.4]
  assign storesToCheck_0_10 = _T_2228 ? _T_7781 : _T_7788; // @[LoadQueue.scala 131:10:@8791.4]
  assign _T_7794 = 4'hb <= offsetQ_0; // @[LoadQueue.scala 131:81:@8794.4]
  assign _T_7795 = _T_6302 & _T_7794; // @[LoadQueue.scala 131:72:@8795.4]
  assign _T_7797 = offsetQ_0 < 4'hb; // @[LoadQueue.scala 132:33:@8796.4]
  assign _T_7800 = _T_7797 & _T_6311; // @[LoadQueue.scala 132:41:@8798.4]
  assign _T_7802 = _T_7800 == 1'h0; // @[LoadQueue.scala 132:9:@8799.4]
  assign storesToCheck_0_11 = _T_2228 ? _T_7795 : _T_7802; // @[LoadQueue.scala 131:10:@8800.4]
  assign _T_7808 = 4'hc <= offsetQ_0; // @[LoadQueue.scala 131:81:@8803.4]
  assign _T_7809 = _T_6319 & _T_7808; // @[LoadQueue.scala 131:72:@8804.4]
  assign _T_7811 = offsetQ_0 < 4'hc; // @[LoadQueue.scala 132:33:@8805.4]
  assign _T_7814 = _T_7811 & _T_6328; // @[LoadQueue.scala 132:41:@8807.4]
  assign _T_7816 = _T_7814 == 1'h0; // @[LoadQueue.scala 132:9:@8808.4]
  assign storesToCheck_0_12 = _T_2228 ? _T_7809 : _T_7816; // @[LoadQueue.scala 131:10:@8809.4]
  assign _T_7822 = 4'hd <= offsetQ_0; // @[LoadQueue.scala 131:81:@8812.4]
  assign _T_7823 = _T_6336 & _T_7822; // @[LoadQueue.scala 131:72:@8813.4]
  assign _T_7825 = offsetQ_0 < 4'hd; // @[LoadQueue.scala 132:33:@8814.4]
  assign _T_7828 = _T_7825 & _T_6345; // @[LoadQueue.scala 132:41:@8816.4]
  assign _T_7830 = _T_7828 == 1'h0; // @[LoadQueue.scala 132:9:@8817.4]
  assign storesToCheck_0_13 = _T_2228 ? _T_7823 : _T_7830; // @[LoadQueue.scala 131:10:@8818.4]
  assign _T_7836 = 4'he <= offsetQ_0; // @[LoadQueue.scala 131:81:@8821.4]
  assign _T_7837 = _T_6353 & _T_7836; // @[LoadQueue.scala 131:72:@8822.4]
  assign _T_7839 = offsetQ_0 < 4'he; // @[LoadQueue.scala 132:33:@8823.4]
  assign _T_7842 = _T_7839 & _T_6362; // @[LoadQueue.scala 132:41:@8825.4]
  assign _T_7844 = _T_7842 == 1'h0; // @[LoadQueue.scala 132:9:@8826.4]
  assign storesToCheck_0_14 = _T_2228 ? _T_7837 : _T_7844; // @[LoadQueue.scala 131:10:@8827.4]
  assign _T_7850 = 4'hf <= offsetQ_0; // @[LoadQueue.scala 131:81:@8830.4]
  assign storesToCheck_0_15 = _T_2228 ? _T_7850 : 1'h1; // @[LoadQueue.scala 131:10:@8836.4]
  assign storesToCheck_1_0 = _T_2258 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@8878.4]
  assign _T_7900 = 4'h1 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8881.4]
  assign _T_7901 = _T_6132 & _T_7900; // @[LoadQueue.scala 131:72:@8882.4]
  assign _T_7903 = offsetQ_1 < 4'h1; // @[LoadQueue.scala 132:33:@8883.4]
  assign _T_7906 = _T_7903 & _T_6141; // @[LoadQueue.scala 132:41:@8885.4]
  assign _T_7908 = _T_7906 == 1'h0; // @[LoadQueue.scala 132:9:@8886.4]
  assign storesToCheck_1_1 = _T_2258 ? _T_7901 : _T_7908; // @[LoadQueue.scala 131:10:@8887.4]
  assign _T_7914 = 4'h2 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8890.4]
  assign _T_7915 = _T_6149 & _T_7914; // @[LoadQueue.scala 131:72:@8891.4]
  assign _T_7917 = offsetQ_1 < 4'h2; // @[LoadQueue.scala 132:33:@8892.4]
  assign _T_7920 = _T_7917 & _T_6158; // @[LoadQueue.scala 132:41:@8894.4]
  assign _T_7922 = _T_7920 == 1'h0; // @[LoadQueue.scala 132:9:@8895.4]
  assign storesToCheck_1_2 = _T_2258 ? _T_7915 : _T_7922; // @[LoadQueue.scala 131:10:@8896.4]
  assign _T_7928 = 4'h3 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8899.4]
  assign _T_7929 = _T_6166 & _T_7928; // @[LoadQueue.scala 131:72:@8900.4]
  assign _T_7931 = offsetQ_1 < 4'h3; // @[LoadQueue.scala 132:33:@8901.4]
  assign _T_7934 = _T_7931 & _T_6175; // @[LoadQueue.scala 132:41:@8903.4]
  assign _T_7936 = _T_7934 == 1'h0; // @[LoadQueue.scala 132:9:@8904.4]
  assign storesToCheck_1_3 = _T_2258 ? _T_7929 : _T_7936; // @[LoadQueue.scala 131:10:@8905.4]
  assign _T_7942 = 4'h4 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8908.4]
  assign _T_7943 = _T_6183 & _T_7942; // @[LoadQueue.scala 131:72:@8909.4]
  assign _T_7945 = offsetQ_1 < 4'h4; // @[LoadQueue.scala 132:33:@8910.4]
  assign _T_7948 = _T_7945 & _T_6192; // @[LoadQueue.scala 132:41:@8912.4]
  assign _T_7950 = _T_7948 == 1'h0; // @[LoadQueue.scala 132:9:@8913.4]
  assign storesToCheck_1_4 = _T_2258 ? _T_7943 : _T_7950; // @[LoadQueue.scala 131:10:@8914.4]
  assign _T_7956 = 4'h5 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8917.4]
  assign _T_7957 = _T_6200 & _T_7956; // @[LoadQueue.scala 131:72:@8918.4]
  assign _T_7959 = offsetQ_1 < 4'h5; // @[LoadQueue.scala 132:33:@8919.4]
  assign _T_7962 = _T_7959 & _T_6209; // @[LoadQueue.scala 132:41:@8921.4]
  assign _T_7964 = _T_7962 == 1'h0; // @[LoadQueue.scala 132:9:@8922.4]
  assign storesToCheck_1_5 = _T_2258 ? _T_7957 : _T_7964; // @[LoadQueue.scala 131:10:@8923.4]
  assign _T_7970 = 4'h6 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8926.4]
  assign _T_7971 = _T_6217 & _T_7970; // @[LoadQueue.scala 131:72:@8927.4]
  assign _T_7973 = offsetQ_1 < 4'h6; // @[LoadQueue.scala 132:33:@8928.4]
  assign _T_7976 = _T_7973 & _T_6226; // @[LoadQueue.scala 132:41:@8930.4]
  assign _T_7978 = _T_7976 == 1'h0; // @[LoadQueue.scala 132:9:@8931.4]
  assign storesToCheck_1_6 = _T_2258 ? _T_7971 : _T_7978; // @[LoadQueue.scala 131:10:@8932.4]
  assign _T_7984 = 4'h7 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8935.4]
  assign _T_7985 = _T_6234 & _T_7984; // @[LoadQueue.scala 131:72:@8936.4]
  assign _T_7987 = offsetQ_1 < 4'h7; // @[LoadQueue.scala 132:33:@8937.4]
  assign _T_7990 = _T_7987 & _T_6243; // @[LoadQueue.scala 132:41:@8939.4]
  assign _T_7992 = _T_7990 == 1'h0; // @[LoadQueue.scala 132:9:@8940.4]
  assign storesToCheck_1_7 = _T_2258 ? _T_7985 : _T_7992; // @[LoadQueue.scala 131:10:@8941.4]
  assign _T_7998 = 4'h8 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8944.4]
  assign _T_7999 = _T_6251 & _T_7998; // @[LoadQueue.scala 131:72:@8945.4]
  assign _T_8001 = offsetQ_1 < 4'h8; // @[LoadQueue.scala 132:33:@8946.4]
  assign _T_8004 = _T_8001 & _T_6260; // @[LoadQueue.scala 132:41:@8948.4]
  assign _T_8006 = _T_8004 == 1'h0; // @[LoadQueue.scala 132:9:@8949.4]
  assign storesToCheck_1_8 = _T_2258 ? _T_7999 : _T_8006; // @[LoadQueue.scala 131:10:@8950.4]
  assign _T_8012 = 4'h9 <= offsetQ_1; // @[LoadQueue.scala 131:81:@8953.4]
  assign _T_8013 = _T_6268 & _T_8012; // @[LoadQueue.scala 131:72:@8954.4]
  assign _T_8015 = offsetQ_1 < 4'h9; // @[LoadQueue.scala 132:33:@8955.4]
  assign _T_8018 = _T_8015 & _T_6277; // @[LoadQueue.scala 132:41:@8957.4]
  assign _T_8020 = _T_8018 == 1'h0; // @[LoadQueue.scala 132:9:@8958.4]
  assign storesToCheck_1_9 = _T_2258 ? _T_8013 : _T_8020; // @[LoadQueue.scala 131:10:@8959.4]
  assign _T_8026 = 4'ha <= offsetQ_1; // @[LoadQueue.scala 131:81:@8962.4]
  assign _T_8027 = _T_6285 & _T_8026; // @[LoadQueue.scala 131:72:@8963.4]
  assign _T_8029 = offsetQ_1 < 4'ha; // @[LoadQueue.scala 132:33:@8964.4]
  assign _T_8032 = _T_8029 & _T_6294; // @[LoadQueue.scala 132:41:@8966.4]
  assign _T_8034 = _T_8032 == 1'h0; // @[LoadQueue.scala 132:9:@8967.4]
  assign storesToCheck_1_10 = _T_2258 ? _T_8027 : _T_8034; // @[LoadQueue.scala 131:10:@8968.4]
  assign _T_8040 = 4'hb <= offsetQ_1; // @[LoadQueue.scala 131:81:@8971.4]
  assign _T_8041 = _T_6302 & _T_8040; // @[LoadQueue.scala 131:72:@8972.4]
  assign _T_8043 = offsetQ_1 < 4'hb; // @[LoadQueue.scala 132:33:@8973.4]
  assign _T_8046 = _T_8043 & _T_6311; // @[LoadQueue.scala 132:41:@8975.4]
  assign _T_8048 = _T_8046 == 1'h0; // @[LoadQueue.scala 132:9:@8976.4]
  assign storesToCheck_1_11 = _T_2258 ? _T_8041 : _T_8048; // @[LoadQueue.scala 131:10:@8977.4]
  assign _T_8054 = 4'hc <= offsetQ_1; // @[LoadQueue.scala 131:81:@8980.4]
  assign _T_8055 = _T_6319 & _T_8054; // @[LoadQueue.scala 131:72:@8981.4]
  assign _T_8057 = offsetQ_1 < 4'hc; // @[LoadQueue.scala 132:33:@8982.4]
  assign _T_8060 = _T_8057 & _T_6328; // @[LoadQueue.scala 132:41:@8984.4]
  assign _T_8062 = _T_8060 == 1'h0; // @[LoadQueue.scala 132:9:@8985.4]
  assign storesToCheck_1_12 = _T_2258 ? _T_8055 : _T_8062; // @[LoadQueue.scala 131:10:@8986.4]
  assign _T_8068 = 4'hd <= offsetQ_1; // @[LoadQueue.scala 131:81:@8989.4]
  assign _T_8069 = _T_6336 & _T_8068; // @[LoadQueue.scala 131:72:@8990.4]
  assign _T_8071 = offsetQ_1 < 4'hd; // @[LoadQueue.scala 132:33:@8991.4]
  assign _T_8074 = _T_8071 & _T_6345; // @[LoadQueue.scala 132:41:@8993.4]
  assign _T_8076 = _T_8074 == 1'h0; // @[LoadQueue.scala 132:9:@8994.4]
  assign storesToCheck_1_13 = _T_2258 ? _T_8069 : _T_8076; // @[LoadQueue.scala 131:10:@8995.4]
  assign _T_8082 = 4'he <= offsetQ_1; // @[LoadQueue.scala 131:81:@8998.4]
  assign _T_8083 = _T_6353 & _T_8082; // @[LoadQueue.scala 131:72:@8999.4]
  assign _T_8085 = offsetQ_1 < 4'he; // @[LoadQueue.scala 132:33:@9000.4]
  assign _T_8088 = _T_8085 & _T_6362; // @[LoadQueue.scala 132:41:@9002.4]
  assign _T_8090 = _T_8088 == 1'h0; // @[LoadQueue.scala 132:9:@9003.4]
  assign storesToCheck_1_14 = _T_2258 ? _T_8083 : _T_8090; // @[LoadQueue.scala 131:10:@9004.4]
  assign _T_8096 = 4'hf <= offsetQ_1; // @[LoadQueue.scala 131:81:@9007.4]
  assign storesToCheck_1_15 = _T_2258 ? _T_8096 : 1'h1; // @[LoadQueue.scala 131:10:@9013.4]
  assign storesToCheck_2_0 = _T_2288 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9055.4]
  assign _T_8146 = 4'h1 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9058.4]
  assign _T_8147 = _T_6132 & _T_8146; // @[LoadQueue.scala 131:72:@9059.4]
  assign _T_8149 = offsetQ_2 < 4'h1; // @[LoadQueue.scala 132:33:@9060.4]
  assign _T_8152 = _T_8149 & _T_6141; // @[LoadQueue.scala 132:41:@9062.4]
  assign _T_8154 = _T_8152 == 1'h0; // @[LoadQueue.scala 132:9:@9063.4]
  assign storesToCheck_2_1 = _T_2288 ? _T_8147 : _T_8154; // @[LoadQueue.scala 131:10:@9064.4]
  assign _T_8160 = 4'h2 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9067.4]
  assign _T_8161 = _T_6149 & _T_8160; // @[LoadQueue.scala 131:72:@9068.4]
  assign _T_8163 = offsetQ_2 < 4'h2; // @[LoadQueue.scala 132:33:@9069.4]
  assign _T_8166 = _T_8163 & _T_6158; // @[LoadQueue.scala 132:41:@9071.4]
  assign _T_8168 = _T_8166 == 1'h0; // @[LoadQueue.scala 132:9:@9072.4]
  assign storesToCheck_2_2 = _T_2288 ? _T_8161 : _T_8168; // @[LoadQueue.scala 131:10:@9073.4]
  assign _T_8174 = 4'h3 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9076.4]
  assign _T_8175 = _T_6166 & _T_8174; // @[LoadQueue.scala 131:72:@9077.4]
  assign _T_8177 = offsetQ_2 < 4'h3; // @[LoadQueue.scala 132:33:@9078.4]
  assign _T_8180 = _T_8177 & _T_6175; // @[LoadQueue.scala 132:41:@9080.4]
  assign _T_8182 = _T_8180 == 1'h0; // @[LoadQueue.scala 132:9:@9081.4]
  assign storesToCheck_2_3 = _T_2288 ? _T_8175 : _T_8182; // @[LoadQueue.scala 131:10:@9082.4]
  assign _T_8188 = 4'h4 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9085.4]
  assign _T_8189 = _T_6183 & _T_8188; // @[LoadQueue.scala 131:72:@9086.4]
  assign _T_8191 = offsetQ_2 < 4'h4; // @[LoadQueue.scala 132:33:@9087.4]
  assign _T_8194 = _T_8191 & _T_6192; // @[LoadQueue.scala 132:41:@9089.4]
  assign _T_8196 = _T_8194 == 1'h0; // @[LoadQueue.scala 132:9:@9090.4]
  assign storesToCheck_2_4 = _T_2288 ? _T_8189 : _T_8196; // @[LoadQueue.scala 131:10:@9091.4]
  assign _T_8202 = 4'h5 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9094.4]
  assign _T_8203 = _T_6200 & _T_8202; // @[LoadQueue.scala 131:72:@9095.4]
  assign _T_8205 = offsetQ_2 < 4'h5; // @[LoadQueue.scala 132:33:@9096.4]
  assign _T_8208 = _T_8205 & _T_6209; // @[LoadQueue.scala 132:41:@9098.4]
  assign _T_8210 = _T_8208 == 1'h0; // @[LoadQueue.scala 132:9:@9099.4]
  assign storesToCheck_2_5 = _T_2288 ? _T_8203 : _T_8210; // @[LoadQueue.scala 131:10:@9100.4]
  assign _T_8216 = 4'h6 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9103.4]
  assign _T_8217 = _T_6217 & _T_8216; // @[LoadQueue.scala 131:72:@9104.4]
  assign _T_8219 = offsetQ_2 < 4'h6; // @[LoadQueue.scala 132:33:@9105.4]
  assign _T_8222 = _T_8219 & _T_6226; // @[LoadQueue.scala 132:41:@9107.4]
  assign _T_8224 = _T_8222 == 1'h0; // @[LoadQueue.scala 132:9:@9108.4]
  assign storesToCheck_2_6 = _T_2288 ? _T_8217 : _T_8224; // @[LoadQueue.scala 131:10:@9109.4]
  assign _T_8230 = 4'h7 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9112.4]
  assign _T_8231 = _T_6234 & _T_8230; // @[LoadQueue.scala 131:72:@9113.4]
  assign _T_8233 = offsetQ_2 < 4'h7; // @[LoadQueue.scala 132:33:@9114.4]
  assign _T_8236 = _T_8233 & _T_6243; // @[LoadQueue.scala 132:41:@9116.4]
  assign _T_8238 = _T_8236 == 1'h0; // @[LoadQueue.scala 132:9:@9117.4]
  assign storesToCheck_2_7 = _T_2288 ? _T_8231 : _T_8238; // @[LoadQueue.scala 131:10:@9118.4]
  assign _T_8244 = 4'h8 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9121.4]
  assign _T_8245 = _T_6251 & _T_8244; // @[LoadQueue.scala 131:72:@9122.4]
  assign _T_8247 = offsetQ_2 < 4'h8; // @[LoadQueue.scala 132:33:@9123.4]
  assign _T_8250 = _T_8247 & _T_6260; // @[LoadQueue.scala 132:41:@9125.4]
  assign _T_8252 = _T_8250 == 1'h0; // @[LoadQueue.scala 132:9:@9126.4]
  assign storesToCheck_2_8 = _T_2288 ? _T_8245 : _T_8252; // @[LoadQueue.scala 131:10:@9127.4]
  assign _T_8258 = 4'h9 <= offsetQ_2; // @[LoadQueue.scala 131:81:@9130.4]
  assign _T_8259 = _T_6268 & _T_8258; // @[LoadQueue.scala 131:72:@9131.4]
  assign _T_8261 = offsetQ_2 < 4'h9; // @[LoadQueue.scala 132:33:@9132.4]
  assign _T_8264 = _T_8261 & _T_6277; // @[LoadQueue.scala 132:41:@9134.4]
  assign _T_8266 = _T_8264 == 1'h0; // @[LoadQueue.scala 132:9:@9135.4]
  assign storesToCheck_2_9 = _T_2288 ? _T_8259 : _T_8266; // @[LoadQueue.scala 131:10:@9136.4]
  assign _T_8272 = 4'ha <= offsetQ_2; // @[LoadQueue.scala 131:81:@9139.4]
  assign _T_8273 = _T_6285 & _T_8272; // @[LoadQueue.scala 131:72:@9140.4]
  assign _T_8275 = offsetQ_2 < 4'ha; // @[LoadQueue.scala 132:33:@9141.4]
  assign _T_8278 = _T_8275 & _T_6294; // @[LoadQueue.scala 132:41:@9143.4]
  assign _T_8280 = _T_8278 == 1'h0; // @[LoadQueue.scala 132:9:@9144.4]
  assign storesToCheck_2_10 = _T_2288 ? _T_8273 : _T_8280; // @[LoadQueue.scala 131:10:@9145.4]
  assign _T_8286 = 4'hb <= offsetQ_2; // @[LoadQueue.scala 131:81:@9148.4]
  assign _T_8287 = _T_6302 & _T_8286; // @[LoadQueue.scala 131:72:@9149.4]
  assign _T_8289 = offsetQ_2 < 4'hb; // @[LoadQueue.scala 132:33:@9150.4]
  assign _T_8292 = _T_8289 & _T_6311; // @[LoadQueue.scala 132:41:@9152.4]
  assign _T_8294 = _T_8292 == 1'h0; // @[LoadQueue.scala 132:9:@9153.4]
  assign storesToCheck_2_11 = _T_2288 ? _T_8287 : _T_8294; // @[LoadQueue.scala 131:10:@9154.4]
  assign _T_8300 = 4'hc <= offsetQ_2; // @[LoadQueue.scala 131:81:@9157.4]
  assign _T_8301 = _T_6319 & _T_8300; // @[LoadQueue.scala 131:72:@9158.4]
  assign _T_8303 = offsetQ_2 < 4'hc; // @[LoadQueue.scala 132:33:@9159.4]
  assign _T_8306 = _T_8303 & _T_6328; // @[LoadQueue.scala 132:41:@9161.4]
  assign _T_8308 = _T_8306 == 1'h0; // @[LoadQueue.scala 132:9:@9162.4]
  assign storesToCheck_2_12 = _T_2288 ? _T_8301 : _T_8308; // @[LoadQueue.scala 131:10:@9163.4]
  assign _T_8314 = 4'hd <= offsetQ_2; // @[LoadQueue.scala 131:81:@9166.4]
  assign _T_8315 = _T_6336 & _T_8314; // @[LoadQueue.scala 131:72:@9167.4]
  assign _T_8317 = offsetQ_2 < 4'hd; // @[LoadQueue.scala 132:33:@9168.4]
  assign _T_8320 = _T_8317 & _T_6345; // @[LoadQueue.scala 132:41:@9170.4]
  assign _T_8322 = _T_8320 == 1'h0; // @[LoadQueue.scala 132:9:@9171.4]
  assign storesToCheck_2_13 = _T_2288 ? _T_8315 : _T_8322; // @[LoadQueue.scala 131:10:@9172.4]
  assign _T_8328 = 4'he <= offsetQ_2; // @[LoadQueue.scala 131:81:@9175.4]
  assign _T_8329 = _T_6353 & _T_8328; // @[LoadQueue.scala 131:72:@9176.4]
  assign _T_8331 = offsetQ_2 < 4'he; // @[LoadQueue.scala 132:33:@9177.4]
  assign _T_8334 = _T_8331 & _T_6362; // @[LoadQueue.scala 132:41:@9179.4]
  assign _T_8336 = _T_8334 == 1'h0; // @[LoadQueue.scala 132:9:@9180.4]
  assign storesToCheck_2_14 = _T_2288 ? _T_8329 : _T_8336; // @[LoadQueue.scala 131:10:@9181.4]
  assign _T_8342 = 4'hf <= offsetQ_2; // @[LoadQueue.scala 131:81:@9184.4]
  assign storesToCheck_2_15 = _T_2288 ? _T_8342 : 1'h1; // @[LoadQueue.scala 131:10:@9190.4]
  assign storesToCheck_3_0 = _T_2318 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9232.4]
  assign _T_8392 = 4'h1 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9235.4]
  assign _T_8393 = _T_6132 & _T_8392; // @[LoadQueue.scala 131:72:@9236.4]
  assign _T_8395 = offsetQ_3 < 4'h1; // @[LoadQueue.scala 132:33:@9237.4]
  assign _T_8398 = _T_8395 & _T_6141; // @[LoadQueue.scala 132:41:@9239.4]
  assign _T_8400 = _T_8398 == 1'h0; // @[LoadQueue.scala 132:9:@9240.4]
  assign storesToCheck_3_1 = _T_2318 ? _T_8393 : _T_8400; // @[LoadQueue.scala 131:10:@9241.4]
  assign _T_8406 = 4'h2 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9244.4]
  assign _T_8407 = _T_6149 & _T_8406; // @[LoadQueue.scala 131:72:@9245.4]
  assign _T_8409 = offsetQ_3 < 4'h2; // @[LoadQueue.scala 132:33:@9246.4]
  assign _T_8412 = _T_8409 & _T_6158; // @[LoadQueue.scala 132:41:@9248.4]
  assign _T_8414 = _T_8412 == 1'h0; // @[LoadQueue.scala 132:9:@9249.4]
  assign storesToCheck_3_2 = _T_2318 ? _T_8407 : _T_8414; // @[LoadQueue.scala 131:10:@9250.4]
  assign _T_8420 = 4'h3 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9253.4]
  assign _T_8421 = _T_6166 & _T_8420; // @[LoadQueue.scala 131:72:@9254.4]
  assign _T_8423 = offsetQ_3 < 4'h3; // @[LoadQueue.scala 132:33:@9255.4]
  assign _T_8426 = _T_8423 & _T_6175; // @[LoadQueue.scala 132:41:@9257.4]
  assign _T_8428 = _T_8426 == 1'h0; // @[LoadQueue.scala 132:9:@9258.4]
  assign storesToCheck_3_3 = _T_2318 ? _T_8421 : _T_8428; // @[LoadQueue.scala 131:10:@9259.4]
  assign _T_8434 = 4'h4 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9262.4]
  assign _T_8435 = _T_6183 & _T_8434; // @[LoadQueue.scala 131:72:@9263.4]
  assign _T_8437 = offsetQ_3 < 4'h4; // @[LoadQueue.scala 132:33:@9264.4]
  assign _T_8440 = _T_8437 & _T_6192; // @[LoadQueue.scala 132:41:@9266.4]
  assign _T_8442 = _T_8440 == 1'h0; // @[LoadQueue.scala 132:9:@9267.4]
  assign storesToCheck_3_4 = _T_2318 ? _T_8435 : _T_8442; // @[LoadQueue.scala 131:10:@9268.4]
  assign _T_8448 = 4'h5 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9271.4]
  assign _T_8449 = _T_6200 & _T_8448; // @[LoadQueue.scala 131:72:@9272.4]
  assign _T_8451 = offsetQ_3 < 4'h5; // @[LoadQueue.scala 132:33:@9273.4]
  assign _T_8454 = _T_8451 & _T_6209; // @[LoadQueue.scala 132:41:@9275.4]
  assign _T_8456 = _T_8454 == 1'h0; // @[LoadQueue.scala 132:9:@9276.4]
  assign storesToCheck_3_5 = _T_2318 ? _T_8449 : _T_8456; // @[LoadQueue.scala 131:10:@9277.4]
  assign _T_8462 = 4'h6 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9280.4]
  assign _T_8463 = _T_6217 & _T_8462; // @[LoadQueue.scala 131:72:@9281.4]
  assign _T_8465 = offsetQ_3 < 4'h6; // @[LoadQueue.scala 132:33:@9282.4]
  assign _T_8468 = _T_8465 & _T_6226; // @[LoadQueue.scala 132:41:@9284.4]
  assign _T_8470 = _T_8468 == 1'h0; // @[LoadQueue.scala 132:9:@9285.4]
  assign storesToCheck_3_6 = _T_2318 ? _T_8463 : _T_8470; // @[LoadQueue.scala 131:10:@9286.4]
  assign _T_8476 = 4'h7 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9289.4]
  assign _T_8477 = _T_6234 & _T_8476; // @[LoadQueue.scala 131:72:@9290.4]
  assign _T_8479 = offsetQ_3 < 4'h7; // @[LoadQueue.scala 132:33:@9291.4]
  assign _T_8482 = _T_8479 & _T_6243; // @[LoadQueue.scala 132:41:@9293.4]
  assign _T_8484 = _T_8482 == 1'h0; // @[LoadQueue.scala 132:9:@9294.4]
  assign storesToCheck_3_7 = _T_2318 ? _T_8477 : _T_8484; // @[LoadQueue.scala 131:10:@9295.4]
  assign _T_8490 = 4'h8 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9298.4]
  assign _T_8491 = _T_6251 & _T_8490; // @[LoadQueue.scala 131:72:@9299.4]
  assign _T_8493 = offsetQ_3 < 4'h8; // @[LoadQueue.scala 132:33:@9300.4]
  assign _T_8496 = _T_8493 & _T_6260; // @[LoadQueue.scala 132:41:@9302.4]
  assign _T_8498 = _T_8496 == 1'h0; // @[LoadQueue.scala 132:9:@9303.4]
  assign storesToCheck_3_8 = _T_2318 ? _T_8491 : _T_8498; // @[LoadQueue.scala 131:10:@9304.4]
  assign _T_8504 = 4'h9 <= offsetQ_3; // @[LoadQueue.scala 131:81:@9307.4]
  assign _T_8505 = _T_6268 & _T_8504; // @[LoadQueue.scala 131:72:@9308.4]
  assign _T_8507 = offsetQ_3 < 4'h9; // @[LoadQueue.scala 132:33:@9309.4]
  assign _T_8510 = _T_8507 & _T_6277; // @[LoadQueue.scala 132:41:@9311.4]
  assign _T_8512 = _T_8510 == 1'h0; // @[LoadQueue.scala 132:9:@9312.4]
  assign storesToCheck_3_9 = _T_2318 ? _T_8505 : _T_8512; // @[LoadQueue.scala 131:10:@9313.4]
  assign _T_8518 = 4'ha <= offsetQ_3; // @[LoadQueue.scala 131:81:@9316.4]
  assign _T_8519 = _T_6285 & _T_8518; // @[LoadQueue.scala 131:72:@9317.4]
  assign _T_8521 = offsetQ_3 < 4'ha; // @[LoadQueue.scala 132:33:@9318.4]
  assign _T_8524 = _T_8521 & _T_6294; // @[LoadQueue.scala 132:41:@9320.4]
  assign _T_8526 = _T_8524 == 1'h0; // @[LoadQueue.scala 132:9:@9321.4]
  assign storesToCheck_3_10 = _T_2318 ? _T_8519 : _T_8526; // @[LoadQueue.scala 131:10:@9322.4]
  assign _T_8532 = 4'hb <= offsetQ_3; // @[LoadQueue.scala 131:81:@9325.4]
  assign _T_8533 = _T_6302 & _T_8532; // @[LoadQueue.scala 131:72:@9326.4]
  assign _T_8535 = offsetQ_3 < 4'hb; // @[LoadQueue.scala 132:33:@9327.4]
  assign _T_8538 = _T_8535 & _T_6311; // @[LoadQueue.scala 132:41:@9329.4]
  assign _T_8540 = _T_8538 == 1'h0; // @[LoadQueue.scala 132:9:@9330.4]
  assign storesToCheck_3_11 = _T_2318 ? _T_8533 : _T_8540; // @[LoadQueue.scala 131:10:@9331.4]
  assign _T_8546 = 4'hc <= offsetQ_3; // @[LoadQueue.scala 131:81:@9334.4]
  assign _T_8547 = _T_6319 & _T_8546; // @[LoadQueue.scala 131:72:@9335.4]
  assign _T_8549 = offsetQ_3 < 4'hc; // @[LoadQueue.scala 132:33:@9336.4]
  assign _T_8552 = _T_8549 & _T_6328; // @[LoadQueue.scala 132:41:@9338.4]
  assign _T_8554 = _T_8552 == 1'h0; // @[LoadQueue.scala 132:9:@9339.4]
  assign storesToCheck_3_12 = _T_2318 ? _T_8547 : _T_8554; // @[LoadQueue.scala 131:10:@9340.4]
  assign _T_8560 = 4'hd <= offsetQ_3; // @[LoadQueue.scala 131:81:@9343.4]
  assign _T_8561 = _T_6336 & _T_8560; // @[LoadQueue.scala 131:72:@9344.4]
  assign _T_8563 = offsetQ_3 < 4'hd; // @[LoadQueue.scala 132:33:@9345.4]
  assign _T_8566 = _T_8563 & _T_6345; // @[LoadQueue.scala 132:41:@9347.4]
  assign _T_8568 = _T_8566 == 1'h0; // @[LoadQueue.scala 132:9:@9348.4]
  assign storesToCheck_3_13 = _T_2318 ? _T_8561 : _T_8568; // @[LoadQueue.scala 131:10:@9349.4]
  assign _T_8574 = 4'he <= offsetQ_3; // @[LoadQueue.scala 131:81:@9352.4]
  assign _T_8575 = _T_6353 & _T_8574; // @[LoadQueue.scala 131:72:@9353.4]
  assign _T_8577 = offsetQ_3 < 4'he; // @[LoadQueue.scala 132:33:@9354.4]
  assign _T_8580 = _T_8577 & _T_6362; // @[LoadQueue.scala 132:41:@9356.4]
  assign _T_8582 = _T_8580 == 1'h0; // @[LoadQueue.scala 132:9:@9357.4]
  assign storesToCheck_3_14 = _T_2318 ? _T_8575 : _T_8582; // @[LoadQueue.scala 131:10:@9358.4]
  assign _T_8588 = 4'hf <= offsetQ_3; // @[LoadQueue.scala 131:81:@9361.4]
  assign storesToCheck_3_15 = _T_2318 ? _T_8588 : 1'h1; // @[LoadQueue.scala 131:10:@9367.4]
  assign storesToCheck_4_0 = _T_2348 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9409.4]
  assign _T_8638 = 4'h1 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9412.4]
  assign _T_8639 = _T_6132 & _T_8638; // @[LoadQueue.scala 131:72:@9413.4]
  assign _T_8641 = offsetQ_4 < 4'h1; // @[LoadQueue.scala 132:33:@9414.4]
  assign _T_8644 = _T_8641 & _T_6141; // @[LoadQueue.scala 132:41:@9416.4]
  assign _T_8646 = _T_8644 == 1'h0; // @[LoadQueue.scala 132:9:@9417.4]
  assign storesToCheck_4_1 = _T_2348 ? _T_8639 : _T_8646; // @[LoadQueue.scala 131:10:@9418.4]
  assign _T_8652 = 4'h2 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9421.4]
  assign _T_8653 = _T_6149 & _T_8652; // @[LoadQueue.scala 131:72:@9422.4]
  assign _T_8655 = offsetQ_4 < 4'h2; // @[LoadQueue.scala 132:33:@9423.4]
  assign _T_8658 = _T_8655 & _T_6158; // @[LoadQueue.scala 132:41:@9425.4]
  assign _T_8660 = _T_8658 == 1'h0; // @[LoadQueue.scala 132:9:@9426.4]
  assign storesToCheck_4_2 = _T_2348 ? _T_8653 : _T_8660; // @[LoadQueue.scala 131:10:@9427.4]
  assign _T_8666 = 4'h3 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9430.4]
  assign _T_8667 = _T_6166 & _T_8666; // @[LoadQueue.scala 131:72:@9431.4]
  assign _T_8669 = offsetQ_4 < 4'h3; // @[LoadQueue.scala 132:33:@9432.4]
  assign _T_8672 = _T_8669 & _T_6175; // @[LoadQueue.scala 132:41:@9434.4]
  assign _T_8674 = _T_8672 == 1'h0; // @[LoadQueue.scala 132:9:@9435.4]
  assign storesToCheck_4_3 = _T_2348 ? _T_8667 : _T_8674; // @[LoadQueue.scala 131:10:@9436.4]
  assign _T_8680 = 4'h4 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9439.4]
  assign _T_8681 = _T_6183 & _T_8680; // @[LoadQueue.scala 131:72:@9440.4]
  assign _T_8683 = offsetQ_4 < 4'h4; // @[LoadQueue.scala 132:33:@9441.4]
  assign _T_8686 = _T_8683 & _T_6192; // @[LoadQueue.scala 132:41:@9443.4]
  assign _T_8688 = _T_8686 == 1'h0; // @[LoadQueue.scala 132:9:@9444.4]
  assign storesToCheck_4_4 = _T_2348 ? _T_8681 : _T_8688; // @[LoadQueue.scala 131:10:@9445.4]
  assign _T_8694 = 4'h5 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9448.4]
  assign _T_8695 = _T_6200 & _T_8694; // @[LoadQueue.scala 131:72:@9449.4]
  assign _T_8697 = offsetQ_4 < 4'h5; // @[LoadQueue.scala 132:33:@9450.4]
  assign _T_8700 = _T_8697 & _T_6209; // @[LoadQueue.scala 132:41:@9452.4]
  assign _T_8702 = _T_8700 == 1'h0; // @[LoadQueue.scala 132:9:@9453.4]
  assign storesToCheck_4_5 = _T_2348 ? _T_8695 : _T_8702; // @[LoadQueue.scala 131:10:@9454.4]
  assign _T_8708 = 4'h6 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9457.4]
  assign _T_8709 = _T_6217 & _T_8708; // @[LoadQueue.scala 131:72:@9458.4]
  assign _T_8711 = offsetQ_4 < 4'h6; // @[LoadQueue.scala 132:33:@9459.4]
  assign _T_8714 = _T_8711 & _T_6226; // @[LoadQueue.scala 132:41:@9461.4]
  assign _T_8716 = _T_8714 == 1'h0; // @[LoadQueue.scala 132:9:@9462.4]
  assign storesToCheck_4_6 = _T_2348 ? _T_8709 : _T_8716; // @[LoadQueue.scala 131:10:@9463.4]
  assign _T_8722 = 4'h7 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9466.4]
  assign _T_8723 = _T_6234 & _T_8722; // @[LoadQueue.scala 131:72:@9467.4]
  assign _T_8725 = offsetQ_4 < 4'h7; // @[LoadQueue.scala 132:33:@9468.4]
  assign _T_8728 = _T_8725 & _T_6243; // @[LoadQueue.scala 132:41:@9470.4]
  assign _T_8730 = _T_8728 == 1'h0; // @[LoadQueue.scala 132:9:@9471.4]
  assign storesToCheck_4_7 = _T_2348 ? _T_8723 : _T_8730; // @[LoadQueue.scala 131:10:@9472.4]
  assign _T_8736 = 4'h8 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9475.4]
  assign _T_8737 = _T_6251 & _T_8736; // @[LoadQueue.scala 131:72:@9476.4]
  assign _T_8739 = offsetQ_4 < 4'h8; // @[LoadQueue.scala 132:33:@9477.4]
  assign _T_8742 = _T_8739 & _T_6260; // @[LoadQueue.scala 132:41:@9479.4]
  assign _T_8744 = _T_8742 == 1'h0; // @[LoadQueue.scala 132:9:@9480.4]
  assign storesToCheck_4_8 = _T_2348 ? _T_8737 : _T_8744; // @[LoadQueue.scala 131:10:@9481.4]
  assign _T_8750 = 4'h9 <= offsetQ_4; // @[LoadQueue.scala 131:81:@9484.4]
  assign _T_8751 = _T_6268 & _T_8750; // @[LoadQueue.scala 131:72:@9485.4]
  assign _T_8753 = offsetQ_4 < 4'h9; // @[LoadQueue.scala 132:33:@9486.4]
  assign _T_8756 = _T_8753 & _T_6277; // @[LoadQueue.scala 132:41:@9488.4]
  assign _T_8758 = _T_8756 == 1'h0; // @[LoadQueue.scala 132:9:@9489.4]
  assign storesToCheck_4_9 = _T_2348 ? _T_8751 : _T_8758; // @[LoadQueue.scala 131:10:@9490.4]
  assign _T_8764 = 4'ha <= offsetQ_4; // @[LoadQueue.scala 131:81:@9493.4]
  assign _T_8765 = _T_6285 & _T_8764; // @[LoadQueue.scala 131:72:@9494.4]
  assign _T_8767 = offsetQ_4 < 4'ha; // @[LoadQueue.scala 132:33:@9495.4]
  assign _T_8770 = _T_8767 & _T_6294; // @[LoadQueue.scala 132:41:@9497.4]
  assign _T_8772 = _T_8770 == 1'h0; // @[LoadQueue.scala 132:9:@9498.4]
  assign storesToCheck_4_10 = _T_2348 ? _T_8765 : _T_8772; // @[LoadQueue.scala 131:10:@9499.4]
  assign _T_8778 = 4'hb <= offsetQ_4; // @[LoadQueue.scala 131:81:@9502.4]
  assign _T_8779 = _T_6302 & _T_8778; // @[LoadQueue.scala 131:72:@9503.4]
  assign _T_8781 = offsetQ_4 < 4'hb; // @[LoadQueue.scala 132:33:@9504.4]
  assign _T_8784 = _T_8781 & _T_6311; // @[LoadQueue.scala 132:41:@9506.4]
  assign _T_8786 = _T_8784 == 1'h0; // @[LoadQueue.scala 132:9:@9507.4]
  assign storesToCheck_4_11 = _T_2348 ? _T_8779 : _T_8786; // @[LoadQueue.scala 131:10:@9508.4]
  assign _T_8792 = 4'hc <= offsetQ_4; // @[LoadQueue.scala 131:81:@9511.4]
  assign _T_8793 = _T_6319 & _T_8792; // @[LoadQueue.scala 131:72:@9512.4]
  assign _T_8795 = offsetQ_4 < 4'hc; // @[LoadQueue.scala 132:33:@9513.4]
  assign _T_8798 = _T_8795 & _T_6328; // @[LoadQueue.scala 132:41:@9515.4]
  assign _T_8800 = _T_8798 == 1'h0; // @[LoadQueue.scala 132:9:@9516.4]
  assign storesToCheck_4_12 = _T_2348 ? _T_8793 : _T_8800; // @[LoadQueue.scala 131:10:@9517.4]
  assign _T_8806 = 4'hd <= offsetQ_4; // @[LoadQueue.scala 131:81:@9520.4]
  assign _T_8807 = _T_6336 & _T_8806; // @[LoadQueue.scala 131:72:@9521.4]
  assign _T_8809 = offsetQ_4 < 4'hd; // @[LoadQueue.scala 132:33:@9522.4]
  assign _T_8812 = _T_8809 & _T_6345; // @[LoadQueue.scala 132:41:@9524.4]
  assign _T_8814 = _T_8812 == 1'h0; // @[LoadQueue.scala 132:9:@9525.4]
  assign storesToCheck_4_13 = _T_2348 ? _T_8807 : _T_8814; // @[LoadQueue.scala 131:10:@9526.4]
  assign _T_8820 = 4'he <= offsetQ_4; // @[LoadQueue.scala 131:81:@9529.4]
  assign _T_8821 = _T_6353 & _T_8820; // @[LoadQueue.scala 131:72:@9530.4]
  assign _T_8823 = offsetQ_4 < 4'he; // @[LoadQueue.scala 132:33:@9531.4]
  assign _T_8826 = _T_8823 & _T_6362; // @[LoadQueue.scala 132:41:@9533.4]
  assign _T_8828 = _T_8826 == 1'h0; // @[LoadQueue.scala 132:9:@9534.4]
  assign storesToCheck_4_14 = _T_2348 ? _T_8821 : _T_8828; // @[LoadQueue.scala 131:10:@9535.4]
  assign _T_8834 = 4'hf <= offsetQ_4; // @[LoadQueue.scala 131:81:@9538.4]
  assign storesToCheck_4_15 = _T_2348 ? _T_8834 : 1'h1; // @[LoadQueue.scala 131:10:@9544.4]
  assign storesToCheck_5_0 = _T_2378 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9586.4]
  assign _T_8884 = 4'h1 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9589.4]
  assign _T_8885 = _T_6132 & _T_8884; // @[LoadQueue.scala 131:72:@9590.4]
  assign _T_8887 = offsetQ_5 < 4'h1; // @[LoadQueue.scala 132:33:@9591.4]
  assign _T_8890 = _T_8887 & _T_6141; // @[LoadQueue.scala 132:41:@9593.4]
  assign _T_8892 = _T_8890 == 1'h0; // @[LoadQueue.scala 132:9:@9594.4]
  assign storesToCheck_5_1 = _T_2378 ? _T_8885 : _T_8892; // @[LoadQueue.scala 131:10:@9595.4]
  assign _T_8898 = 4'h2 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9598.4]
  assign _T_8899 = _T_6149 & _T_8898; // @[LoadQueue.scala 131:72:@9599.4]
  assign _T_8901 = offsetQ_5 < 4'h2; // @[LoadQueue.scala 132:33:@9600.4]
  assign _T_8904 = _T_8901 & _T_6158; // @[LoadQueue.scala 132:41:@9602.4]
  assign _T_8906 = _T_8904 == 1'h0; // @[LoadQueue.scala 132:9:@9603.4]
  assign storesToCheck_5_2 = _T_2378 ? _T_8899 : _T_8906; // @[LoadQueue.scala 131:10:@9604.4]
  assign _T_8912 = 4'h3 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9607.4]
  assign _T_8913 = _T_6166 & _T_8912; // @[LoadQueue.scala 131:72:@9608.4]
  assign _T_8915 = offsetQ_5 < 4'h3; // @[LoadQueue.scala 132:33:@9609.4]
  assign _T_8918 = _T_8915 & _T_6175; // @[LoadQueue.scala 132:41:@9611.4]
  assign _T_8920 = _T_8918 == 1'h0; // @[LoadQueue.scala 132:9:@9612.4]
  assign storesToCheck_5_3 = _T_2378 ? _T_8913 : _T_8920; // @[LoadQueue.scala 131:10:@9613.4]
  assign _T_8926 = 4'h4 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9616.4]
  assign _T_8927 = _T_6183 & _T_8926; // @[LoadQueue.scala 131:72:@9617.4]
  assign _T_8929 = offsetQ_5 < 4'h4; // @[LoadQueue.scala 132:33:@9618.4]
  assign _T_8932 = _T_8929 & _T_6192; // @[LoadQueue.scala 132:41:@9620.4]
  assign _T_8934 = _T_8932 == 1'h0; // @[LoadQueue.scala 132:9:@9621.4]
  assign storesToCheck_5_4 = _T_2378 ? _T_8927 : _T_8934; // @[LoadQueue.scala 131:10:@9622.4]
  assign _T_8940 = 4'h5 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9625.4]
  assign _T_8941 = _T_6200 & _T_8940; // @[LoadQueue.scala 131:72:@9626.4]
  assign _T_8943 = offsetQ_5 < 4'h5; // @[LoadQueue.scala 132:33:@9627.4]
  assign _T_8946 = _T_8943 & _T_6209; // @[LoadQueue.scala 132:41:@9629.4]
  assign _T_8948 = _T_8946 == 1'h0; // @[LoadQueue.scala 132:9:@9630.4]
  assign storesToCheck_5_5 = _T_2378 ? _T_8941 : _T_8948; // @[LoadQueue.scala 131:10:@9631.4]
  assign _T_8954 = 4'h6 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9634.4]
  assign _T_8955 = _T_6217 & _T_8954; // @[LoadQueue.scala 131:72:@9635.4]
  assign _T_8957 = offsetQ_5 < 4'h6; // @[LoadQueue.scala 132:33:@9636.4]
  assign _T_8960 = _T_8957 & _T_6226; // @[LoadQueue.scala 132:41:@9638.4]
  assign _T_8962 = _T_8960 == 1'h0; // @[LoadQueue.scala 132:9:@9639.4]
  assign storesToCheck_5_6 = _T_2378 ? _T_8955 : _T_8962; // @[LoadQueue.scala 131:10:@9640.4]
  assign _T_8968 = 4'h7 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9643.4]
  assign _T_8969 = _T_6234 & _T_8968; // @[LoadQueue.scala 131:72:@9644.4]
  assign _T_8971 = offsetQ_5 < 4'h7; // @[LoadQueue.scala 132:33:@9645.4]
  assign _T_8974 = _T_8971 & _T_6243; // @[LoadQueue.scala 132:41:@9647.4]
  assign _T_8976 = _T_8974 == 1'h0; // @[LoadQueue.scala 132:9:@9648.4]
  assign storesToCheck_5_7 = _T_2378 ? _T_8969 : _T_8976; // @[LoadQueue.scala 131:10:@9649.4]
  assign _T_8982 = 4'h8 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9652.4]
  assign _T_8983 = _T_6251 & _T_8982; // @[LoadQueue.scala 131:72:@9653.4]
  assign _T_8985 = offsetQ_5 < 4'h8; // @[LoadQueue.scala 132:33:@9654.4]
  assign _T_8988 = _T_8985 & _T_6260; // @[LoadQueue.scala 132:41:@9656.4]
  assign _T_8990 = _T_8988 == 1'h0; // @[LoadQueue.scala 132:9:@9657.4]
  assign storesToCheck_5_8 = _T_2378 ? _T_8983 : _T_8990; // @[LoadQueue.scala 131:10:@9658.4]
  assign _T_8996 = 4'h9 <= offsetQ_5; // @[LoadQueue.scala 131:81:@9661.4]
  assign _T_8997 = _T_6268 & _T_8996; // @[LoadQueue.scala 131:72:@9662.4]
  assign _T_8999 = offsetQ_5 < 4'h9; // @[LoadQueue.scala 132:33:@9663.4]
  assign _T_9002 = _T_8999 & _T_6277; // @[LoadQueue.scala 132:41:@9665.4]
  assign _T_9004 = _T_9002 == 1'h0; // @[LoadQueue.scala 132:9:@9666.4]
  assign storesToCheck_5_9 = _T_2378 ? _T_8997 : _T_9004; // @[LoadQueue.scala 131:10:@9667.4]
  assign _T_9010 = 4'ha <= offsetQ_5; // @[LoadQueue.scala 131:81:@9670.4]
  assign _T_9011 = _T_6285 & _T_9010; // @[LoadQueue.scala 131:72:@9671.4]
  assign _T_9013 = offsetQ_5 < 4'ha; // @[LoadQueue.scala 132:33:@9672.4]
  assign _T_9016 = _T_9013 & _T_6294; // @[LoadQueue.scala 132:41:@9674.4]
  assign _T_9018 = _T_9016 == 1'h0; // @[LoadQueue.scala 132:9:@9675.4]
  assign storesToCheck_5_10 = _T_2378 ? _T_9011 : _T_9018; // @[LoadQueue.scala 131:10:@9676.4]
  assign _T_9024 = 4'hb <= offsetQ_5; // @[LoadQueue.scala 131:81:@9679.4]
  assign _T_9025 = _T_6302 & _T_9024; // @[LoadQueue.scala 131:72:@9680.4]
  assign _T_9027 = offsetQ_5 < 4'hb; // @[LoadQueue.scala 132:33:@9681.4]
  assign _T_9030 = _T_9027 & _T_6311; // @[LoadQueue.scala 132:41:@9683.4]
  assign _T_9032 = _T_9030 == 1'h0; // @[LoadQueue.scala 132:9:@9684.4]
  assign storesToCheck_5_11 = _T_2378 ? _T_9025 : _T_9032; // @[LoadQueue.scala 131:10:@9685.4]
  assign _T_9038 = 4'hc <= offsetQ_5; // @[LoadQueue.scala 131:81:@9688.4]
  assign _T_9039 = _T_6319 & _T_9038; // @[LoadQueue.scala 131:72:@9689.4]
  assign _T_9041 = offsetQ_5 < 4'hc; // @[LoadQueue.scala 132:33:@9690.4]
  assign _T_9044 = _T_9041 & _T_6328; // @[LoadQueue.scala 132:41:@9692.4]
  assign _T_9046 = _T_9044 == 1'h0; // @[LoadQueue.scala 132:9:@9693.4]
  assign storesToCheck_5_12 = _T_2378 ? _T_9039 : _T_9046; // @[LoadQueue.scala 131:10:@9694.4]
  assign _T_9052 = 4'hd <= offsetQ_5; // @[LoadQueue.scala 131:81:@9697.4]
  assign _T_9053 = _T_6336 & _T_9052; // @[LoadQueue.scala 131:72:@9698.4]
  assign _T_9055 = offsetQ_5 < 4'hd; // @[LoadQueue.scala 132:33:@9699.4]
  assign _T_9058 = _T_9055 & _T_6345; // @[LoadQueue.scala 132:41:@9701.4]
  assign _T_9060 = _T_9058 == 1'h0; // @[LoadQueue.scala 132:9:@9702.4]
  assign storesToCheck_5_13 = _T_2378 ? _T_9053 : _T_9060; // @[LoadQueue.scala 131:10:@9703.4]
  assign _T_9066 = 4'he <= offsetQ_5; // @[LoadQueue.scala 131:81:@9706.4]
  assign _T_9067 = _T_6353 & _T_9066; // @[LoadQueue.scala 131:72:@9707.4]
  assign _T_9069 = offsetQ_5 < 4'he; // @[LoadQueue.scala 132:33:@9708.4]
  assign _T_9072 = _T_9069 & _T_6362; // @[LoadQueue.scala 132:41:@9710.4]
  assign _T_9074 = _T_9072 == 1'h0; // @[LoadQueue.scala 132:9:@9711.4]
  assign storesToCheck_5_14 = _T_2378 ? _T_9067 : _T_9074; // @[LoadQueue.scala 131:10:@9712.4]
  assign _T_9080 = 4'hf <= offsetQ_5; // @[LoadQueue.scala 131:81:@9715.4]
  assign storesToCheck_5_15 = _T_2378 ? _T_9080 : 1'h1; // @[LoadQueue.scala 131:10:@9721.4]
  assign storesToCheck_6_0 = _T_2408 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9763.4]
  assign _T_9130 = 4'h1 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9766.4]
  assign _T_9131 = _T_6132 & _T_9130; // @[LoadQueue.scala 131:72:@9767.4]
  assign _T_9133 = offsetQ_6 < 4'h1; // @[LoadQueue.scala 132:33:@9768.4]
  assign _T_9136 = _T_9133 & _T_6141; // @[LoadQueue.scala 132:41:@9770.4]
  assign _T_9138 = _T_9136 == 1'h0; // @[LoadQueue.scala 132:9:@9771.4]
  assign storesToCheck_6_1 = _T_2408 ? _T_9131 : _T_9138; // @[LoadQueue.scala 131:10:@9772.4]
  assign _T_9144 = 4'h2 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9775.4]
  assign _T_9145 = _T_6149 & _T_9144; // @[LoadQueue.scala 131:72:@9776.4]
  assign _T_9147 = offsetQ_6 < 4'h2; // @[LoadQueue.scala 132:33:@9777.4]
  assign _T_9150 = _T_9147 & _T_6158; // @[LoadQueue.scala 132:41:@9779.4]
  assign _T_9152 = _T_9150 == 1'h0; // @[LoadQueue.scala 132:9:@9780.4]
  assign storesToCheck_6_2 = _T_2408 ? _T_9145 : _T_9152; // @[LoadQueue.scala 131:10:@9781.4]
  assign _T_9158 = 4'h3 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9784.4]
  assign _T_9159 = _T_6166 & _T_9158; // @[LoadQueue.scala 131:72:@9785.4]
  assign _T_9161 = offsetQ_6 < 4'h3; // @[LoadQueue.scala 132:33:@9786.4]
  assign _T_9164 = _T_9161 & _T_6175; // @[LoadQueue.scala 132:41:@9788.4]
  assign _T_9166 = _T_9164 == 1'h0; // @[LoadQueue.scala 132:9:@9789.4]
  assign storesToCheck_6_3 = _T_2408 ? _T_9159 : _T_9166; // @[LoadQueue.scala 131:10:@9790.4]
  assign _T_9172 = 4'h4 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9793.4]
  assign _T_9173 = _T_6183 & _T_9172; // @[LoadQueue.scala 131:72:@9794.4]
  assign _T_9175 = offsetQ_6 < 4'h4; // @[LoadQueue.scala 132:33:@9795.4]
  assign _T_9178 = _T_9175 & _T_6192; // @[LoadQueue.scala 132:41:@9797.4]
  assign _T_9180 = _T_9178 == 1'h0; // @[LoadQueue.scala 132:9:@9798.4]
  assign storesToCheck_6_4 = _T_2408 ? _T_9173 : _T_9180; // @[LoadQueue.scala 131:10:@9799.4]
  assign _T_9186 = 4'h5 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9802.4]
  assign _T_9187 = _T_6200 & _T_9186; // @[LoadQueue.scala 131:72:@9803.4]
  assign _T_9189 = offsetQ_6 < 4'h5; // @[LoadQueue.scala 132:33:@9804.4]
  assign _T_9192 = _T_9189 & _T_6209; // @[LoadQueue.scala 132:41:@9806.4]
  assign _T_9194 = _T_9192 == 1'h0; // @[LoadQueue.scala 132:9:@9807.4]
  assign storesToCheck_6_5 = _T_2408 ? _T_9187 : _T_9194; // @[LoadQueue.scala 131:10:@9808.4]
  assign _T_9200 = 4'h6 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9811.4]
  assign _T_9201 = _T_6217 & _T_9200; // @[LoadQueue.scala 131:72:@9812.4]
  assign _T_9203 = offsetQ_6 < 4'h6; // @[LoadQueue.scala 132:33:@9813.4]
  assign _T_9206 = _T_9203 & _T_6226; // @[LoadQueue.scala 132:41:@9815.4]
  assign _T_9208 = _T_9206 == 1'h0; // @[LoadQueue.scala 132:9:@9816.4]
  assign storesToCheck_6_6 = _T_2408 ? _T_9201 : _T_9208; // @[LoadQueue.scala 131:10:@9817.4]
  assign _T_9214 = 4'h7 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9820.4]
  assign _T_9215 = _T_6234 & _T_9214; // @[LoadQueue.scala 131:72:@9821.4]
  assign _T_9217 = offsetQ_6 < 4'h7; // @[LoadQueue.scala 132:33:@9822.4]
  assign _T_9220 = _T_9217 & _T_6243; // @[LoadQueue.scala 132:41:@9824.4]
  assign _T_9222 = _T_9220 == 1'h0; // @[LoadQueue.scala 132:9:@9825.4]
  assign storesToCheck_6_7 = _T_2408 ? _T_9215 : _T_9222; // @[LoadQueue.scala 131:10:@9826.4]
  assign _T_9228 = 4'h8 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9829.4]
  assign _T_9229 = _T_6251 & _T_9228; // @[LoadQueue.scala 131:72:@9830.4]
  assign _T_9231 = offsetQ_6 < 4'h8; // @[LoadQueue.scala 132:33:@9831.4]
  assign _T_9234 = _T_9231 & _T_6260; // @[LoadQueue.scala 132:41:@9833.4]
  assign _T_9236 = _T_9234 == 1'h0; // @[LoadQueue.scala 132:9:@9834.4]
  assign storesToCheck_6_8 = _T_2408 ? _T_9229 : _T_9236; // @[LoadQueue.scala 131:10:@9835.4]
  assign _T_9242 = 4'h9 <= offsetQ_6; // @[LoadQueue.scala 131:81:@9838.4]
  assign _T_9243 = _T_6268 & _T_9242; // @[LoadQueue.scala 131:72:@9839.4]
  assign _T_9245 = offsetQ_6 < 4'h9; // @[LoadQueue.scala 132:33:@9840.4]
  assign _T_9248 = _T_9245 & _T_6277; // @[LoadQueue.scala 132:41:@9842.4]
  assign _T_9250 = _T_9248 == 1'h0; // @[LoadQueue.scala 132:9:@9843.4]
  assign storesToCheck_6_9 = _T_2408 ? _T_9243 : _T_9250; // @[LoadQueue.scala 131:10:@9844.4]
  assign _T_9256 = 4'ha <= offsetQ_6; // @[LoadQueue.scala 131:81:@9847.4]
  assign _T_9257 = _T_6285 & _T_9256; // @[LoadQueue.scala 131:72:@9848.4]
  assign _T_9259 = offsetQ_6 < 4'ha; // @[LoadQueue.scala 132:33:@9849.4]
  assign _T_9262 = _T_9259 & _T_6294; // @[LoadQueue.scala 132:41:@9851.4]
  assign _T_9264 = _T_9262 == 1'h0; // @[LoadQueue.scala 132:9:@9852.4]
  assign storesToCheck_6_10 = _T_2408 ? _T_9257 : _T_9264; // @[LoadQueue.scala 131:10:@9853.4]
  assign _T_9270 = 4'hb <= offsetQ_6; // @[LoadQueue.scala 131:81:@9856.4]
  assign _T_9271 = _T_6302 & _T_9270; // @[LoadQueue.scala 131:72:@9857.4]
  assign _T_9273 = offsetQ_6 < 4'hb; // @[LoadQueue.scala 132:33:@9858.4]
  assign _T_9276 = _T_9273 & _T_6311; // @[LoadQueue.scala 132:41:@9860.4]
  assign _T_9278 = _T_9276 == 1'h0; // @[LoadQueue.scala 132:9:@9861.4]
  assign storesToCheck_6_11 = _T_2408 ? _T_9271 : _T_9278; // @[LoadQueue.scala 131:10:@9862.4]
  assign _T_9284 = 4'hc <= offsetQ_6; // @[LoadQueue.scala 131:81:@9865.4]
  assign _T_9285 = _T_6319 & _T_9284; // @[LoadQueue.scala 131:72:@9866.4]
  assign _T_9287 = offsetQ_6 < 4'hc; // @[LoadQueue.scala 132:33:@9867.4]
  assign _T_9290 = _T_9287 & _T_6328; // @[LoadQueue.scala 132:41:@9869.4]
  assign _T_9292 = _T_9290 == 1'h0; // @[LoadQueue.scala 132:9:@9870.4]
  assign storesToCheck_6_12 = _T_2408 ? _T_9285 : _T_9292; // @[LoadQueue.scala 131:10:@9871.4]
  assign _T_9298 = 4'hd <= offsetQ_6; // @[LoadQueue.scala 131:81:@9874.4]
  assign _T_9299 = _T_6336 & _T_9298; // @[LoadQueue.scala 131:72:@9875.4]
  assign _T_9301 = offsetQ_6 < 4'hd; // @[LoadQueue.scala 132:33:@9876.4]
  assign _T_9304 = _T_9301 & _T_6345; // @[LoadQueue.scala 132:41:@9878.4]
  assign _T_9306 = _T_9304 == 1'h0; // @[LoadQueue.scala 132:9:@9879.4]
  assign storesToCheck_6_13 = _T_2408 ? _T_9299 : _T_9306; // @[LoadQueue.scala 131:10:@9880.4]
  assign _T_9312 = 4'he <= offsetQ_6; // @[LoadQueue.scala 131:81:@9883.4]
  assign _T_9313 = _T_6353 & _T_9312; // @[LoadQueue.scala 131:72:@9884.4]
  assign _T_9315 = offsetQ_6 < 4'he; // @[LoadQueue.scala 132:33:@9885.4]
  assign _T_9318 = _T_9315 & _T_6362; // @[LoadQueue.scala 132:41:@9887.4]
  assign _T_9320 = _T_9318 == 1'h0; // @[LoadQueue.scala 132:9:@9888.4]
  assign storesToCheck_6_14 = _T_2408 ? _T_9313 : _T_9320; // @[LoadQueue.scala 131:10:@9889.4]
  assign _T_9326 = 4'hf <= offsetQ_6; // @[LoadQueue.scala 131:81:@9892.4]
  assign storesToCheck_6_15 = _T_2408 ? _T_9326 : 1'h1; // @[LoadQueue.scala 131:10:@9898.4]
  assign storesToCheck_7_0 = _T_2438 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@9940.4]
  assign _T_9376 = 4'h1 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9943.4]
  assign _T_9377 = _T_6132 & _T_9376; // @[LoadQueue.scala 131:72:@9944.4]
  assign _T_9379 = offsetQ_7 < 4'h1; // @[LoadQueue.scala 132:33:@9945.4]
  assign _T_9382 = _T_9379 & _T_6141; // @[LoadQueue.scala 132:41:@9947.4]
  assign _T_9384 = _T_9382 == 1'h0; // @[LoadQueue.scala 132:9:@9948.4]
  assign storesToCheck_7_1 = _T_2438 ? _T_9377 : _T_9384; // @[LoadQueue.scala 131:10:@9949.4]
  assign _T_9390 = 4'h2 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9952.4]
  assign _T_9391 = _T_6149 & _T_9390; // @[LoadQueue.scala 131:72:@9953.4]
  assign _T_9393 = offsetQ_7 < 4'h2; // @[LoadQueue.scala 132:33:@9954.4]
  assign _T_9396 = _T_9393 & _T_6158; // @[LoadQueue.scala 132:41:@9956.4]
  assign _T_9398 = _T_9396 == 1'h0; // @[LoadQueue.scala 132:9:@9957.4]
  assign storesToCheck_7_2 = _T_2438 ? _T_9391 : _T_9398; // @[LoadQueue.scala 131:10:@9958.4]
  assign _T_9404 = 4'h3 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9961.4]
  assign _T_9405 = _T_6166 & _T_9404; // @[LoadQueue.scala 131:72:@9962.4]
  assign _T_9407 = offsetQ_7 < 4'h3; // @[LoadQueue.scala 132:33:@9963.4]
  assign _T_9410 = _T_9407 & _T_6175; // @[LoadQueue.scala 132:41:@9965.4]
  assign _T_9412 = _T_9410 == 1'h0; // @[LoadQueue.scala 132:9:@9966.4]
  assign storesToCheck_7_3 = _T_2438 ? _T_9405 : _T_9412; // @[LoadQueue.scala 131:10:@9967.4]
  assign _T_9418 = 4'h4 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9970.4]
  assign _T_9419 = _T_6183 & _T_9418; // @[LoadQueue.scala 131:72:@9971.4]
  assign _T_9421 = offsetQ_7 < 4'h4; // @[LoadQueue.scala 132:33:@9972.4]
  assign _T_9424 = _T_9421 & _T_6192; // @[LoadQueue.scala 132:41:@9974.4]
  assign _T_9426 = _T_9424 == 1'h0; // @[LoadQueue.scala 132:9:@9975.4]
  assign storesToCheck_7_4 = _T_2438 ? _T_9419 : _T_9426; // @[LoadQueue.scala 131:10:@9976.4]
  assign _T_9432 = 4'h5 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9979.4]
  assign _T_9433 = _T_6200 & _T_9432; // @[LoadQueue.scala 131:72:@9980.4]
  assign _T_9435 = offsetQ_7 < 4'h5; // @[LoadQueue.scala 132:33:@9981.4]
  assign _T_9438 = _T_9435 & _T_6209; // @[LoadQueue.scala 132:41:@9983.4]
  assign _T_9440 = _T_9438 == 1'h0; // @[LoadQueue.scala 132:9:@9984.4]
  assign storesToCheck_7_5 = _T_2438 ? _T_9433 : _T_9440; // @[LoadQueue.scala 131:10:@9985.4]
  assign _T_9446 = 4'h6 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9988.4]
  assign _T_9447 = _T_6217 & _T_9446; // @[LoadQueue.scala 131:72:@9989.4]
  assign _T_9449 = offsetQ_7 < 4'h6; // @[LoadQueue.scala 132:33:@9990.4]
  assign _T_9452 = _T_9449 & _T_6226; // @[LoadQueue.scala 132:41:@9992.4]
  assign _T_9454 = _T_9452 == 1'h0; // @[LoadQueue.scala 132:9:@9993.4]
  assign storesToCheck_7_6 = _T_2438 ? _T_9447 : _T_9454; // @[LoadQueue.scala 131:10:@9994.4]
  assign _T_9460 = 4'h7 <= offsetQ_7; // @[LoadQueue.scala 131:81:@9997.4]
  assign _T_9461 = _T_6234 & _T_9460; // @[LoadQueue.scala 131:72:@9998.4]
  assign _T_9463 = offsetQ_7 < 4'h7; // @[LoadQueue.scala 132:33:@9999.4]
  assign _T_9466 = _T_9463 & _T_6243; // @[LoadQueue.scala 132:41:@10001.4]
  assign _T_9468 = _T_9466 == 1'h0; // @[LoadQueue.scala 132:9:@10002.4]
  assign storesToCheck_7_7 = _T_2438 ? _T_9461 : _T_9468; // @[LoadQueue.scala 131:10:@10003.4]
  assign _T_9474 = 4'h8 <= offsetQ_7; // @[LoadQueue.scala 131:81:@10006.4]
  assign _T_9475 = _T_6251 & _T_9474; // @[LoadQueue.scala 131:72:@10007.4]
  assign _T_9477 = offsetQ_7 < 4'h8; // @[LoadQueue.scala 132:33:@10008.4]
  assign _T_9480 = _T_9477 & _T_6260; // @[LoadQueue.scala 132:41:@10010.4]
  assign _T_9482 = _T_9480 == 1'h0; // @[LoadQueue.scala 132:9:@10011.4]
  assign storesToCheck_7_8 = _T_2438 ? _T_9475 : _T_9482; // @[LoadQueue.scala 131:10:@10012.4]
  assign _T_9488 = 4'h9 <= offsetQ_7; // @[LoadQueue.scala 131:81:@10015.4]
  assign _T_9489 = _T_6268 & _T_9488; // @[LoadQueue.scala 131:72:@10016.4]
  assign _T_9491 = offsetQ_7 < 4'h9; // @[LoadQueue.scala 132:33:@10017.4]
  assign _T_9494 = _T_9491 & _T_6277; // @[LoadQueue.scala 132:41:@10019.4]
  assign _T_9496 = _T_9494 == 1'h0; // @[LoadQueue.scala 132:9:@10020.4]
  assign storesToCheck_7_9 = _T_2438 ? _T_9489 : _T_9496; // @[LoadQueue.scala 131:10:@10021.4]
  assign _T_9502 = 4'ha <= offsetQ_7; // @[LoadQueue.scala 131:81:@10024.4]
  assign _T_9503 = _T_6285 & _T_9502; // @[LoadQueue.scala 131:72:@10025.4]
  assign _T_9505 = offsetQ_7 < 4'ha; // @[LoadQueue.scala 132:33:@10026.4]
  assign _T_9508 = _T_9505 & _T_6294; // @[LoadQueue.scala 132:41:@10028.4]
  assign _T_9510 = _T_9508 == 1'h0; // @[LoadQueue.scala 132:9:@10029.4]
  assign storesToCheck_7_10 = _T_2438 ? _T_9503 : _T_9510; // @[LoadQueue.scala 131:10:@10030.4]
  assign _T_9516 = 4'hb <= offsetQ_7; // @[LoadQueue.scala 131:81:@10033.4]
  assign _T_9517 = _T_6302 & _T_9516; // @[LoadQueue.scala 131:72:@10034.4]
  assign _T_9519 = offsetQ_7 < 4'hb; // @[LoadQueue.scala 132:33:@10035.4]
  assign _T_9522 = _T_9519 & _T_6311; // @[LoadQueue.scala 132:41:@10037.4]
  assign _T_9524 = _T_9522 == 1'h0; // @[LoadQueue.scala 132:9:@10038.4]
  assign storesToCheck_7_11 = _T_2438 ? _T_9517 : _T_9524; // @[LoadQueue.scala 131:10:@10039.4]
  assign _T_9530 = 4'hc <= offsetQ_7; // @[LoadQueue.scala 131:81:@10042.4]
  assign _T_9531 = _T_6319 & _T_9530; // @[LoadQueue.scala 131:72:@10043.4]
  assign _T_9533 = offsetQ_7 < 4'hc; // @[LoadQueue.scala 132:33:@10044.4]
  assign _T_9536 = _T_9533 & _T_6328; // @[LoadQueue.scala 132:41:@10046.4]
  assign _T_9538 = _T_9536 == 1'h0; // @[LoadQueue.scala 132:9:@10047.4]
  assign storesToCheck_7_12 = _T_2438 ? _T_9531 : _T_9538; // @[LoadQueue.scala 131:10:@10048.4]
  assign _T_9544 = 4'hd <= offsetQ_7; // @[LoadQueue.scala 131:81:@10051.4]
  assign _T_9545 = _T_6336 & _T_9544; // @[LoadQueue.scala 131:72:@10052.4]
  assign _T_9547 = offsetQ_7 < 4'hd; // @[LoadQueue.scala 132:33:@10053.4]
  assign _T_9550 = _T_9547 & _T_6345; // @[LoadQueue.scala 132:41:@10055.4]
  assign _T_9552 = _T_9550 == 1'h0; // @[LoadQueue.scala 132:9:@10056.4]
  assign storesToCheck_7_13 = _T_2438 ? _T_9545 : _T_9552; // @[LoadQueue.scala 131:10:@10057.4]
  assign _T_9558 = 4'he <= offsetQ_7; // @[LoadQueue.scala 131:81:@10060.4]
  assign _T_9559 = _T_6353 & _T_9558; // @[LoadQueue.scala 131:72:@10061.4]
  assign _T_9561 = offsetQ_7 < 4'he; // @[LoadQueue.scala 132:33:@10062.4]
  assign _T_9564 = _T_9561 & _T_6362; // @[LoadQueue.scala 132:41:@10064.4]
  assign _T_9566 = _T_9564 == 1'h0; // @[LoadQueue.scala 132:9:@10065.4]
  assign storesToCheck_7_14 = _T_2438 ? _T_9559 : _T_9566; // @[LoadQueue.scala 131:10:@10066.4]
  assign _T_9572 = 4'hf <= offsetQ_7; // @[LoadQueue.scala 131:81:@10069.4]
  assign storesToCheck_7_15 = _T_2438 ? _T_9572 : 1'h1; // @[LoadQueue.scala 131:10:@10075.4]
  assign storesToCheck_8_0 = _T_2468 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@10117.4]
  assign _T_9622 = 4'h1 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10120.4]
  assign _T_9623 = _T_6132 & _T_9622; // @[LoadQueue.scala 131:72:@10121.4]
  assign _T_9625 = offsetQ_8 < 4'h1; // @[LoadQueue.scala 132:33:@10122.4]
  assign _T_9628 = _T_9625 & _T_6141; // @[LoadQueue.scala 132:41:@10124.4]
  assign _T_9630 = _T_9628 == 1'h0; // @[LoadQueue.scala 132:9:@10125.4]
  assign storesToCheck_8_1 = _T_2468 ? _T_9623 : _T_9630; // @[LoadQueue.scala 131:10:@10126.4]
  assign _T_9636 = 4'h2 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10129.4]
  assign _T_9637 = _T_6149 & _T_9636; // @[LoadQueue.scala 131:72:@10130.4]
  assign _T_9639 = offsetQ_8 < 4'h2; // @[LoadQueue.scala 132:33:@10131.4]
  assign _T_9642 = _T_9639 & _T_6158; // @[LoadQueue.scala 132:41:@10133.4]
  assign _T_9644 = _T_9642 == 1'h0; // @[LoadQueue.scala 132:9:@10134.4]
  assign storesToCheck_8_2 = _T_2468 ? _T_9637 : _T_9644; // @[LoadQueue.scala 131:10:@10135.4]
  assign _T_9650 = 4'h3 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10138.4]
  assign _T_9651 = _T_6166 & _T_9650; // @[LoadQueue.scala 131:72:@10139.4]
  assign _T_9653 = offsetQ_8 < 4'h3; // @[LoadQueue.scala 132:33:@10140.4]
  assign _T_9656 = _T_9653 & _T_6175; // @[LoadQueue.scala 132:41:@10142.4]
  assign _T_9658 = _T_9656 == 1'h0; // @[LoadQueue.scala 132:9:@10143.4]
  assign storesToCheck_8_3 = _T_2468 ? _T_9651 : _T_9658; // @[LoadQueue.scala 131:10:@10144.4]
  assign _T_9664 = 4'h4 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10147.4]
  assign _T_9665 = _T_6183 & _T_9664; // @[LoadQueue.scala 131:72:@10148.4]
  assign _T_9667 = offsetQ_8 < 4'h4; // @[LoadQueue.scala 132:33:@10149.4]
  assign _T_9670 = _T_9667 & _T_6192; // @[LoadQueue.scala 132:41:@10151.4]
  assign _T_9672 = _T_9670 == 1'h0; // @[LoadQueue.scala 132:9:@10152.4]
  assign storesToCheck_8_4 = _T_2468 ? _T_9665 : _T_9672; // @[LoadQueue.scala 131:10:@10153.4]
  assign _T_9678 = 4'h5 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10156.4]
  assign _T_9679 = _T_6200 & _T_9678; // @[LoadQueue.scala 131:72:@10157.4]
  assign _T_9681 = offsetQ_8 < 4'h5; // @[LoadQueue.scala 132:33:@10158.4]
  assign _T_9684 = _T_9681 & _T_6209; // @[LoadQueue.scala 132:41:@10160.4]
  assign _T_9686 = _T_9684 == 1'h0; // @[LoadQueue.scala 132:9:@10161.4]
  assign storesToCheck_8_5 = _T_2468 ? _T_9679 : _T_9686; // @[LoadQueue.scala 131:10:@10162.4]
  assign _T_9692 = 4'h6 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10165.4]
  assign _T_9693 = _T_6217 & _T_9692; // @[LoadQueue.scala 131:72:@10166.4]
  assign _T_9695 = offsetQ_8 < 4'h6; // @[LoadQueue.scala 132:33:@10167.4]
  assign _T_9698 = _T_9695 & _T_6226; // @[LoadQueue.scala 132:41:@10169.4]
  assign _T_9700 = _T_9698 == 1'h0; // @[LoadQueue.scala 132:9:@10170.4]
  assign storesToCheck_8_6 = _T_2468 ? _T_9693 : _T_9700; // @[LoadQueue.scala 131:10:@10171.4]
  assign _T_9706 = 4'h7 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10174.4]
  assign _T_9707 = _T_6234 & _T_9706; // @[LoadQueue.scala 131:72:@10175.4]
  assign _T_9709 = offsetQ_8 < 4'h7; // @[LoadQueue.scala 132:33:@10176.4]
  assign _T_9712 = _T_9709 & _T_6243; // @[LoadQueue.scala 132:41:@10178.4]
  assign _T_9714 = _T_9712 == 1'h0; // @[LoadQueue.scala 132:9:@10179.4]
  assign storesToCheck_8_7 = _T_2468 ? _T_9707 : _T_9714; // @[LoadQueue.scala 131:10:@10180.4]
  assign _T_9720 = 4'h8 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10183.4]
  assign _T_9721 = _T_6251 & _T_9720; // @[LoadQueue.scala 131:72:@10184.4]
  assign _T_9723 = offsetQ_8 < 4'h8; // @[LoadQueue.scala 132:33:@10185.4]
  assign _T_9726 = _T_9723 & _T_6260; // @[LoadQueue.scala 132:41:@10187.4]
  assign _T_9728 = _T_9726 == 1'h0; // @[LoadQueue.scala 132:9:@10188.4]
  assign storesToCheck_8_8 = _T_2468 ? _T_9721 : _T_9728; // @[LoadQueue.scala 131:10:@10189.4]
  assign _T_9734 = 4'h9 <= offsetQ_8; // @[LoadQueue.scala 131:81:@10192.4]
  assign _T_9735 = _T_6268 & _T_9734; // @[LoadQueue.scala 131:72:@10193.4]
  assign _T_9737 = offsetQ_8 < 4'h9; // @[LoadQueue.scala 132:33:@10194.4]
  assign _T_9740 = _T_9737 & _T_6277; // @[LoadQueue.scala 132:41:@10196.4]
  assign _T_9742 = _T_9740 == 1'h0; // @[LoadQueue.scala 132:9:@10197.4]
  assign storesToCheck_8_9 = _T_2468 ? _T_9735 : _T_9742; // @[LoadQueue.scala 131:10:@10198.4]
  assign _T_9748 = 4'ha <= offsetQ_8; // @[LoadQueue.scala 131:81:@10201.4]
  assign _T_9749 = _T_6285 & _T_9748; // @[LoadQueue.scala 131:72:@10202.4]
  assign _T_9751 = offsetQ_8 < 4'ha; // @[LoadQueue.scala 132:33:@10203.4]
  assign _T_9754 = _T_9751 & _T_6294; // @[LoadQueue.scala 132:41:@10205.4]
  assign _T_9756 = _T_9754 == 1'h0; // @[LoadQueue.scala 132:9:@10206.4]
  assign storesToCheck_8_10 = _T_2468 ? _T_9749 : _T_9756; // @[LoadQueue.scala 131:10:@10207.4]
  assign _T_9762 = 4'hb <= offsetQ_8; // @[LoadQueue.scala 131:81:@10210.4]
  assign _T_9763 = _T_6302 & _T_9762; // @[LoadQueue.scala 131:72:@10211.4]
  assign _T_9765 = offsetQ_8 < 4'hb; // @[LoadQueue.scala 132:33:@10212.4]
  assign _T_9768 = _T_9765 & _T_6311; // @[LoadQueue.scala 132:41:@10214.4]
  assign _T_9770 = _T_9768 == 1'h0; // @[LoadQueue.scala 132:9:@10215.4]
  assign storesToCheck_8_11 = _T_2468 ? _T_9763 : _T_9770; // @[LoadQueue.scala 131:10:@10216.4]
  assign _T_9776 = 4'hc <= offsetQ_8; // @[LoadQueue.scala 131:81:@10219.4]
  assign _T_9777 = _T_6319 & _T_9776; // @[LoadQueue.scala 131:72:@10220.4]
  assign _T_9779 = offsetQ_8 < 4'hc; // @[LoadQueue.scala 132:33:@10221.4]
  assign _T_9782 = _T_9779 & _T_6328; // @[LoadQueue.scala 132:41:@10223.4]
  assign _T_9784 = _T_9782 == 1'h0; // @[LoadQueue.scala 132:9:@10224.4]
  assign storesToCheck_8_12 = _T_2468 ? _T_9777 : _T_9784; // @[LoadQueue.scala 131:10:@10225.4]
  assign _T_9790 = 4'hd <= offsetQ_8; // @[LoadQueue.scala 131:81:@10228.4]
  assign _T_9791 = _T_6336 & _T_9790; // @[LoadQueue.scala 131:72:@10229.4]
  assign _T_9793 = offsetQ_8 < 4'hd; // @[LoadQueue.scala 132:33:@10230.4]
  assign _T_9796 = _T_9793 & _T_6345; // @[LoadQueue.scala 132:41:@10232.4]
  assign _T_9798 = _T_9796 == 1'h0; // @[LoadQueue.scala 132:9:@10233.4]
  assign storesToCheck_8_13 = _T_2468 ? _T_9791 : _T_9798; // @[LoadQueue.scala 131:10:@10234.4]
  assign _T_9804 = 4'he <= offsetQ_8; // @[LoadQueue.scala 131:81:@10237.4]
  assign _T_9805 = _T_6353 & _T_9804; // @[LoadQueue.scala 131:72:@10238.4]
  assign _T_9807 = offsetQ_8 < 4'he; // @[LoadQueue.scala 132:33:@10239.4]
  assign _T_9810 = _T_9807 & _T_6362; // @[LoadQueue.scala 132:41:@10241.4]
  assign _T_9812 = _T_9810 == 1'h0; // @[LoadQueue.scala 132:9:@10242.4]
  assign storesToCheck_8_14 = _T_2468 ? _T_9805 : _T_9812; // @[LoadQueue.scala 131:10:@10243.4]
  assign _T_9818 = 4'hf <= offsetQ_8; // @[LoadQueue.scala 131:81:@10246.4]
  assign storesToCheck_8_15 = _T_2468 ? _T_9818 : 1'h1; // @[LoadQueue.scala 131:10:@10252.4]
  assign storesToCheck_9_0 = _T_2498 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@10294.4]
  assign _T_9868 = 4'h1 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10297.4]
  assign _T_9869 = _T_6132 & _T_9868; // @[LoadQueue.scala 131:72:@10298.4]
  assign _T_9871 = offsetQ_9 < 4'h1; // @[LoadQueue.scala 132:33:@10299.4]
  assign _T_9874 = _T_9871 & _T_6141; // @[LoadQueue.scala 132:41:@10301.4]
  assign _T_9876 = _T_9874 == 1'h0; // @[LoadQueue.scala 132:9:@10302.4]
  assign storesToCheck_9_1 = _T_2498 ? _T_9869 : _T_9876; // @[LoadQueue.scala 131:10:@10303.4]
  assign _T_9882 = 4'h2 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10306.4]
  assign _T_9883 = _T_6149 & _T_9882; // @[LoadQueue.scala 131:72:@10307.4]
  assign _T_9885 = offsetQ_9 < 4'h2; // @[LoadQueue.scala 132:33:@10308.4]
  assign _T_9888 = _T_9885 & _T_6158; // @[LoadQueue.scala 132:41:@10310.4]
  assign _T_9890 = _T_9888 == 1'h0; // @[LoadQueue.scala 132:9:@10311.4]
  assign storesToCheck_9_2 = _T_2498 ? _T_9883 : _T_9890; // @[LoadQueue.scala 131:10:@10312.4]
  assign _T_9896 = 4'h3 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10315.4]
  assign _T_9897 = _T_6166 & _T_9896; // @[LoadQueue.scala 131:72:@10316.4]
  assign _T_9899 = offsetQ_9 < 4'h3; // @[LoadQueue.scala 132:33:@10317.4]
  assign _T_9902 = _T_9899 & _T_6175; // @[LoadQueue.scala 132:41:@10319.4]
  assign _T_9904 = _T_9902 == 1'h0; // @[LoadQueue.scala 132:9:@10320.4]
  assign storesToCheck_9_3 = _T_2498 ? _T_9897 : _T_9904; // @[LoadQueue.scala 131:10:@10321.4]
  assign _T_9910 = 4'h4 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10324.4]
  assign _T_9911 = _T_6183 & _T_9910; // @[LoadQueue.scala 131:72:@10325.4]
  assign _T_9913 = offsetQ_9 < 4'h4; // @[LoadQueue.scala 132:33:@10326.4]
  assign _T_9916 = _T_9913 & _T_6192; // @[LoadQueue.scala 132:41:@10328.4]
  assign _T_9918 = _T_9916 == 1'h0; // @[LoadQueue.scala 132:9:@10329.4]
  assign storesToCheck_9_4 = _T_2498 ? _T_9911 : _T_9918; // @[LoadQueue.scala 131:10:@10330.4]
  assign _T_9924 = 4'h5 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10333.4]
  assign _T_9925 = _T_6200 & _T_9924; // @[LoadQueue.scala 131:72:@10334.4]
  assign _T_9927 = offsetQ_9 < 4'h5; // @[LoadQueue.scala 132:33:@10335.4]
  assign _T_9930 = _T_9927 & _T_6209; // @[LoadQueue.scala 132:41:@10337.4]
  assign _T_9932 = _T_9930 == 1'h0; // @[LoadQueue.scala 132:9:@10338.4]
  assign storesToCheck_9_5 = _T_2498 ? _T_9925 : _T_9932; // @[LoadQueue.scala 131:10:@10339.4]
  assign _T_9938 = 4'h6 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10342.4]
  assign _T_9939 = _T_6217 & _T_9938; // @[LoadQueue.scala 131:72:@10343.4]
  assign _T_9941 = offsetQ_9 < 4'h6; // @[LoadQueue.scala 132:33:@10344.4]
  assign _T_9944 = _T_9941 & _T_6226; // @[LoadQueue.scala 132:41:@10346.4]
  assign _T_9946 = _T_9944 == 1'h0; // @[LoadQueue.scala 132:9:@10347.4]
  assign storesToCheck_9_6 = _T_2498 ? _T_9939 : _T_9946; // @[LoadQueue.scala 131:10:@10348.4]
  assign _T_9952 = 4'h7 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10351.4]
  assign _T_9953 = _T_6234 & _T_9952; // @[LoadQueue.scala 131:72:@10352.4]
  assign _T_9955 = offsetQ_9 < 4'h7; // @[LoadQueue.scala 132:33:@10353.4]
  assign _T_9958 = _T_9955 & _T_6243; // @[LoadQueue.scala 132:41:@10355.4]
  assign _T_9960 = _T_9958 == 1'h0; // @[LoadQueue.scala 132:9:@10356.4]
  assign storesToCheck_9_7 = _T_2498 ? _T_9953 : _T_9960; // @[LoadQueue.scala 131:10:@10357.4]
  assign _T_9966 = 4'h8 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10360.4]
  assign _T_9967 = _T_6251 & _T_9966; // @[LoadQueue.scala 131:72:@10361.4]
  assign _T_9969 = offsetQ_9 < 4'h8; // @[LoadQueue.scala 132:33:@10362.4]
  assign _T_9972 = _T_9969 & _T_6260; // @[LoadQueue.scala 132:41:@10364.4]
  assign _T_9974 = _T_9972 == 1'h0; // @[LoadQueue.scala 132:9:@10365.4]
  assign storesToCheck_9_8 = _T_2498 ? _T_9967 : _T_9974; // @[LoadQueue.scala 131:10:@10366.4]
  assign _T_9980 = 4'h9 <= offsetQ_9; // @[LoadQueue.scala 131:81:@10369.4]
  assign _T_9981 = _T_6268 & _T_9980; // @[LoadQueue.scala 131:72:@10370.4]
  assign _T_9983 = offsetQ_9 < 4'h9; // @[LoadQueue.scala 132:33:@10371.4]
  assign _T_9986 = _T_9983 & _T_6277; // @[LoadQueue.scala 132:41:@10373.4]
  assign _T_9988 = _T_9986 == 1'h0; // @[LoadQueue.scala 132:9:@10374.4]
  assign storesToCheck_9_9 = _T_2498 ? _T_9981 : _T_9988; // @[LoadQueue.scala 131:10:@10375.4]
  assign _T_9994 = 4'ha <= offsetQ_9; // @[LoadQueue.scala 131:81:@10378.4]
  assign _T_9995 = _T_6285 & _T_9994; // @[LoadQueue.scala 131:72:@10379.4]
  assign _T_9997 = offsetQ_9 < 4'ha; // @[LoadQueue.scala 132:33:@10380.4]
  assign _T_10000 = _T_9997 & _T_6294; // @[LoadQueue.scala 132:41:@10382.4]
  assign _T_10002 = _T_10000 == 1'h0; // @[LoadQueue.scala 132:9:@10383.4]
  assign storesToCheck_9_10 = _T_2498 ? _T_9995 : _T_10002; // @[LoadQueue.scala 131:10:@10384.4]
  assign _T_10008 = 4'hb <= offsetQ_9; // @[LoadQueue.scala 131:81:@10387.4]
  assign _T_10009 = _T_6302 & _T_10008; // @[LoadQueue.scala 131:72:@10388.4]
  assign _T_10011 = offsetQ_9 < 4'hb; // @[LoadQueue.scala 132:33:@10389.4]
  assign _T_10014 = _T_10011 & _T_6311; // @[LoadQueue.scala 132:41:@10391.4]
  assign _T_10016 = _T_10014 == 1'h0; // @[LoadQueue.scala 132:9:@10392.4]
  assign storesToCheck_9_11 = _T_2498 ? _T_10009 : _T_10016; // @[LoadQueue.scala 131:10:@10393.4]
  assign _T_10022 = 4'hc <= offsetQ_9; // @[LoadQueue.scala 131:81:@10396.4]
  assign _T_10023 = _T_6319 & _T_10022; // @[LoadQueue.scala 131:72:@10397.4]
  assign _T_10025 = offsetQ_9 < 4'hc; // @[LoadQueue.scala 132:33:@10398.4]
  assign _T_10028 = _T_10025 & _T_6328; // @[LoadQueue.scala 132:41:@10400.4]
  assign _T_10030 = _T_10028 == 1'h0; // @[LoadQueue.scala 132:9:@10401.4]
  assign storesToCheck_9_12 = _T_2498 ? _T_10023 : _T_10030; // @[LoadQueue.scala 131:10:@10402.4]
  assign _T_10036 = 4'hd <= offsetQ_9; // @[LoadQueue.scala 131:81:@10405.4]
  assign _T_10037 = _T_6336 & _T_10036; // @[LoadQueue.scala 131:72:@10406.4]
  assign _T_10039 = offsetQ_9 < 4'hd; // @[LoadQueue.scala 132:33:@10407.4]
  assign _T_10042 = _T_10039 & _T_6345; // @[LoadQueue.scala 132:41:@10409.4]
  assign _T_10044 = _T_10042 == 1'h0; // @[LoadQueue.scala 132:9:@10410.4]
  assign storesToCheck_9_13 = _T_2498 ? _T_10037 : _T_10044; // @[LoadQueue.scala 131:10:@10411.4]
  assign _T_10050 = 4'he <= offsetQ_9; // @[LoadQueue.scala 131:81:@10414.4]
  assign _T_10051 = _T_6353 & _T_10050; // @[LoadQueue.scala 131:72:@10415.4]
  assign _T_10053 = offsetQ_9 < 4'he; // @[LoadQueue.scala 132:33:@10416.4]
  assign _T_10056 = _T_10053 & _T_6362; // @[LoadQueue.scala 132:41:@10418.4]
  assign _T_10058 = _T_10056 == 1'h0; // @[LoadQueue.scala 132:9:@10419.4]
  assign storesToCheck_9_14 = _T_2498 ? _T_10051 : _T_10058; // @[LoadQueue.scala 131:10:@10420.4]
  assign _T_10064 = 4'hf <= offsetQ_9; // @[LoadQueue.scala 131:81:@10423.4]
  assign storesToCheck_9_15 = _T_2498 ? _T_10064 : 1'h1; // @[LoadQueue.scala 131:10:@10429.4]
  assign storesToCheck_10_0 = _T_2528 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@10471.4]
  assign _T_10114 = 4'h1 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10474.4]
  assign _T_10115 = _T_6132 & _T_10114; // @[LoadQueue.scala 131:72:@10475.4]
  assign _T_10117 = offsetQ_10 < 4'h1; // @[LoadQueue.scala 132:33:@10476.4]
  assign _T_10120 = _T_10117 & _T_6141; // @[LoadQueue.scala 132:41:@10478.4]
  assign _T_10122 = _T_10120 == 1'h0; // @[LoadQueue.scala 132:9:@10479.4]
  assign storesToCheck_10_1 = _T_2528 ? _T_10115 : _T_10122; // @[LoadQueue.scala 131:10:@10480.4]
  assign _T_10128 = 4'h2 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10483.4]
  assign _T_10129 = _T_6149 & _T_10128; // @[LoadQueue.scala 131:72:@10484.4]
  assign _T_10131 = offsetQ_10 < 4'h2; // @[LoadQueue.scala 132:33:@10485.4]
  assign _T_10134 = _T_10131 & _T_6158; // @[LoadQueue.scala 132:41:@10487.4]
  assign _T_10136 = _T_10134 == 1'h0; // @[LoadQueue.scala 132:9:@10488.4]
  assign storesToCheck_10_2 = _T_2528 ? _T_10129 : _T_10136; // @[LoadQueue.scala 131:10:@10489.4]
  assign _T_10142 = 4'h3 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10492.4]
  assign _T_10143 = _T_6166 & _T_10142; // @[LoadQueue.scala 131:72:@10493.4]
  assign _T_10145 = offsetQ_10 < 4'h3; // @[LoadQueue.scala 132:33:@10494.4]
  assign _T_10148 = _T_10145 & _T_6175; // @[LoadQueue.scala 132:41:@10496.4]
  assign _T_10150 = _T_10148 == 1'h0; // @[LoadQueue.scala 132:9:@10497.4]
  assign storesToCheck_10_3 = _T_2528 ? _T_10143 : _T_10150; // @[LoadQueue.scala 131:10:@10498.4]
  assign _T_10156 = 4'h4 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10501.4]
  assign _T_10157 = _T_6183 & _T_10156; // @[LoadQueue.scala 131:72:@10502.4]
  assign _T_10159 = offsetQ_10 < 4'h4; // @[LoadQueue.scala 132:33:@10503.4]
  assign _T_10162 = _T_10159 & _T_6192; // @[LoadQueue.scala 132:41:@10505.4]
  assign _T_10164 = _T_10162 == 1'h0; // @[LoadQueue.scala 132:9:@10506.4]
  assign storesToCheck_10_4 = _T_2528 ? _T_10157 : _T_10164; // @[LoadQueue.scala 131:10:@10507.4]
  assign _T_10170 = 4'h5 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10510.4]
  assign _T_10171 = _T_6200 & _T_10170; // @[LoadQueue.scala 131:72:@10511.4]
  assign _T_10173 = offsetQ_10 < 4'h5; // @[LoadQueue.scala 132:33:@10512.4]
  assign _T_10176 = _T_10173 & _T_6209; // @[LoadQueue.scala 132:41:@10514.4]
  assign _T_10178 = _T_10176 == 1'h0; // @[LoadQueue.scala 132:9:@10515.4]
  assign storesToCheck_10_5 = _T_2528 ? _T_10171 : _T_10178; // @[LoadQueue.scala 131:10:@10516.4]
  assign _T_10184 = 4'h6 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10519.4]
  assign _T_10185 = _T_6217 & _T_10184; // @[LoadQueue.scala 131:72:@10520.4]
  assign _T_10187 = offsetQ_10 < 4'h6; // @[LoadQueue.scala 132:33:@10521.4]
  assign _T_10190 = _T_10187 & _T_6226; // @[LoadQueue.scala 132:41:@10523.4]
  assign _T_10192 = _T_10190 == 1'h0; // @[LoadQueue.scala 132:9:@10524.4]
  assign storesToCheck_10_6 = _T_2528 ? _T_10185 : _T_10192; // @[LoadQueue.scala 131:10:@10525.4]
  assign _T_10198 = 4'h7 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10528.4]
  assign _T_10199 = _T_6234 & _T_10198; // @[LoadQueue.scala 131:72:@10529.4]
  assign _T_10201 = offsetQ_10 < 4'h7; // @[LoadQueue.scala 132:33:@10530.4]
  assign _T_10204 = _T_10201 & _T_6243; // @[LoadQueue.scala 132:41:@10532.4]
  assign _T_10206 = _T_10204 == 1'h0; // @[LoadQueue.scala 132:9:@10533.4]
  assign storesToCheck_10_7 = _T_2528 ? _T_10199 : _T_10206; // @[LoadQueue.scala 131:10:@10534.4]
  assign _T_10212 = 4'h8 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10537.4]
  assign _T_10213 = _T_6251 & _T_10212; // @[LoadQueue.scala 131:72:@10538.4]
  assign _T_10215 = offsetQ_10 < 4'h8; // @[LoadQueue.scala 132:33:@10539.4]
  assign _T_10218 = _T_10215 & _T_6260; // @[LoadQueue.scala 132:41:@10541.4]
  assign _T_10220 = _T_10218 == 1'h0; // @[LoadQueue.scala 132:9:@10542.4]
  assign storesToCheck_10_8 = _T_2528 ? _T_10213 : _T_10220; // @[LoadQueue.scala 131:10:@10543.4]
  assign _T_10226 = 4'h9 <= offsetQ_10; // @[LoadQueue.scala 131:81:@10546.4]
  assign _T_10227 = _T_6268 & _T_10226; // @[LoadQueue.scala 131:72:@10547.4]
  assign _T_10229 = offsetQ_10 < 4'h9; // @[LoadQueue.scala 132:33:@10548.4]
  assign _T_10232 = _T_10229 & _T_6277; // @[LoadQueue.scala 132:41:@10550.4]
  assign _T_10234 = _T_10232 == 1'h0; // @[LoadQueue.scala 132:9:@10551.4]
  assign storesToCheck_10_9 = _T_2528 ? _T_10227 : _T_10234; // @[LoadQueue.scala 131:10:@10552.4]
  assign _T_10240 = 4'ha <= offsetQ_10; // @[LoadQueue.scala 131:81:@10555.4]
  assign _T_10241 = _T_6285 & _T_10240; // @[LoadQueue.scala 131:72:@10556.4]
  assign _T_10243 = offsetQ_10 < 4'ha; // @[LoadQueue.scala 132:33:@10557.4]
  assign _T_10246 = _T_10243 & _T_6294; // @[LoadQueue.scala 132:41:@10559.4]
  assign _T_10248 = _T_10246 == 1'h0; // @[LoadQueue.scala 132:9:@10560.4]
  assign storesToCheck_10_10 = _T_2528 ? _T_10241 : _T_10248; // @[LoadQueue.scala 131:10:@10561.4]
  assign _T_10254 = 4'hb <= offsetQ_10; // @[LoadQueue.scala 131:81:@10564.4]
  assign _T_10255 = _T_6302 & _T_10254; // @[LoadQueue.scala 131:72:@10565.4]
  assign _T_10257 = offsetQ_10 < 4'hb; // @[LoadQueue.scala 132:33:@10566.4]
  assign _T_10260 = _T_10257 & _T_6311; // @[LoadQueue.scala 132:41:@10568.4]
  assign _T_10262 = _T_10260 == 1'h0; // @[LoadQueue.scala 132:9:@10569.4]
  assign storesToCheck_10_11 = _T_2528 ? _T_10255 : _T_10262; // @[LoadQueue.scala 131:10:@10570.4]
  assign _T_10268 = 4'hc <= offsetQ_10; // @[LoadQueue.scala 131:81:@10573.4]
  assign _T_10269 = _T_6319 & _T_10268; // @[LoadQueue.scala 131:72:@10574.4]
  assign _T_10271 = offsetQ_10 < 4'hc; // @[LoadQueue.scala 132:33:@10575.4]
  assign _T_10274 = _T_10271 & _T_6328; // @[LoadQueue.scala 132:41:@10577.4]
  assign _T_10276 = _T_10274 == 1'h0; // @[LoadQueue.scala 132:9:@10578.4]
  assign storesToCheck_10_12 = _T_2528 ? _T_10269 : _T_10276; // @[LoadQueue.scala 131:10:@10579.4]
  assign _T_10282 = 4'hd <= offsetQ_10; // @[LoadQueue.scala 131:81:@10582.4]
  assign _T_10283 = _T_6336 & _T_10282; // @[LoadQueue.scala 131:72:@10583.4]
  assign _T_10285 = offsetQ_10 < 4'hd; // @[LoadQueue.scala 132:33:@10584.4]
  assign _T_10288 = _T_10285 & _T_6345; // @[LoadQueue.scala 132:41:@10586.4]
  assign _T_10290 = _T_10288 == 1'h0; // @[LoadQueue.scala 132:9:@10587.4]
  assign storesToCheck_10_13 = _T_2528 ? _T_10283 : _T_10290; // @[LoadQueue.scala 131:10:@10588.4]
  assign _T_10296 = 4'he <= offsetQ_10; // @[LoadQueue.scala 131:81:@10591.4]
  assign _T_10297 = _T_6353 & _T_10296; // @[LoadQueue.scala 131:72:@10592.4]
  assign _T_10299 = offsetQ_10 < 4'he; // @[LoadQueue.scala 132:33:@10593.4]
  assign _T_10302 = _T_10299 & _T_6362; // @[LoadQueue.scala 132:41:@10595.4]
  assign _T_10304 = _T_10302 == 1'h0; // @[LoadQueue.scala 132:9:@10596.4]
  assign storesToCheck_10_14 = _T_2528 ? _T_10297 : _T_10304; // @[LoadQueue.scala 131:10:@10597.4]
  assign _T_10310 = 4'hf <= offsetQ_10; // @[LoadQueue.scala 131:81:@10600.4]
  assign storesToCheck_10_15 = _T_2528 ? _T_10310 : 1'h1; // @[LoadQueue.scala 131:10:@10606.4]
  assign storesToCheck_11_0 = _T_2558 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@10648.4]
  assign _T_10360 = 4'h1 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10651.4]
  assign _T_10361 = _T_6132 & _T_10360; // @[LoadQueue.scala 131:72:@10652.4]
  assign _T_10363 = offsetQ_11 < 4'h1; // @[LoadQueue.scala 132:33:@10653.4]
  assign _T_10366 = _T_10363 & _T_6141; // @[LoadQueue.scala 132:41:@10655.4]
  assign _T_10368 = _T_10366 == 1'h0; // @[LoadQueue.scala 132:9:@10656.4]
  assign storesToCheck_11_1 = _T_2558 ? _T_10361 : _T_10368; // @[LoadQueue.scala 131:10:@10657.4]
  assign _T_10374 = 4'h2 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10660.4]
  assign _T_10375 = _T_6149 & _T_10374; // @[LoadQueue.scala 131:72:@10661.4]
  assign _T_10377 = offsetQ_11 < 4'h2; // @[LoadQueue.scala 132:33:@10662.4]
  assign _T_10380 = _T_10377 & _T_6158; // @[LoadQueue.scala 132:41:@10664.4]
  assign _T_10382 = _T_10380 == 1'h0; // @[LoadQueue.scala 132:9:@10665.4]
  assign storesToCheck_11_2 = _T_2558 ? _T_10375 : _T_10382; // @[LoadQueue.scala 131:10:@10666.4]
  assign _T_10388 = 4'h3 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10669.4]
  assign _T_10389 = _T_6166 & _T_10388; // @[LoadQueue.scala 131:72:@10670.4]
  assign _T_10391 = offsetQ_11 < 4'h3; // @[LoadQueue.scala 132:33:@10671.4]
  assign _T_10394 = _T_10391 & _T_6175; // @[LoadQueue.scala 132:41:@10673.4]
  assign _T_10396 = _T_10394 == 1'h0; // @[LoadQueue.scala 132:9:@10674.4]
  assign storesToCheck_11_3 = _T_2558 ? _T_10389 : _T_10396; // @[LoadQueue.scala 131:10:@10675.4]
  assign _T_10402 = 4'h4 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10678.4]
  assign _T_10403 = _T_6183 & _T_10402; // @[LoadQueue.scala 131:72:@10679.4]
  assign _T_10405 = offsetQ_11 < 4'h4; // @[LoadQueue.scala 132:33:@10680.4]
  assign _T_10408 = _T_10405 & _T_6192; // @[LoadQueue.scala 132:41:@10682.4]
  assign _T_10410 = _T_10408 == 1'h0; // @[LoadQueue.scala 132:9:@10683.4]
  assign storesToCheck_11_4 = _T_2558 ? _T_10403 : _T_10410; // @[LoadQueue.scala 131:10:@10684.4]
  assign _T_10416 = 4'h5 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10687.4]
  assign _T_10417 = _T_6200 & _T_10416; // @[LoadQueue.scala 131:72:@10688.4]
  assign _T_10419 = offsetQ_11 < 4'h5; // @[LoadQueue.scala 132:33:@10689.4]
  assign _T_10422 = _T_10419 & _T_6209; // @[LoadQueue.scala 132:41:@10691.4]
  assign _T_10424 = _T_10422 == 1'h0; // @[LoadQueue.scala 132:9:@10692.4]
  assign storesToCheck_11_5 = _T_2558 ? _T_10417 : _T_10424; // @[LoadQueue.scala 131:10:@10693.4]
  assign _T_10430 = 4'h6 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10696.4]
  assign _T_10431 = _T_6217 & _T_10430; // @[LoadQueue.scala 131:72:@10697.4]
  assign _T_10433 = offsetQ_11 < 4'h6; // @[LoadQueue.scala 132:33:@10698.4]
  assign _T_10436 = _T_10433 & _T_6226; // @[LoadQueue.scala 132:41:@10700.4]
  assign _T_10438 = _T_10436 == 1'h0; // @[LoadQueue.scala 132:9:@10701.4]
  assign storesToCheck_11_6 = _T_2558 ? _T_10431 : _T_10438; // @[LoadQueue.scala 131:10:@10702.4]
  assign _T_10444 = 4'h7 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10705.4]
  assign _T_10445 = _T_6234 & _T_10444; // @[LoadQueue.scala 131:72:@10706.4]
  assign _T_10447 = offsetQ_11 < 4'h7; // @[LoadQueue.scala 132:33:@10707.4]
  assign _T_10450 = _T_10447 & _T_6243; // @[LoadQueue.scala 132:41:@10709.4]
  assign _T_10452 = _T_10450 == 1'h0; // @[LoadQueue.scala 132:9:@10710.4]
  assign storesToCheck_11_7 = _T_2558 ? _T_10445 : _T_10452; // @[LoadQueue.scala 131:10:@10711.4]
  assign _T_10458 = 4'h8 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10714.4]
  assign _T_10459 = _T_6251 & _T_10458; // @[LoadQueue.scala 131:72:@10715.4]
  assign _T_10461 = offsetQ_11 < 4'h8; // @[LoadQueue.scala 132:33:@10716.4]
  assign _T_10464 = _T_10461 & _T_6260; // @[LoadQueue.scala 132:41:@10718.4]
  assign _T_10466 = _T_10464 == 1'h0; // @[LoadQueue.scala 132:9:@10719.4]
  assign storesToCheck_11_8 = _T_2558 ? _T_10459 : _T_10466; // @[LoadQueue.scala 131:10:@10720.4]
  assign _T_10472 = 4'h9 <= offsetQ_11; // @[LoadQueue.scala 131:81:@10723.4]
  assign _T_10473 = _T_6268 & _T_10472; // @[LoadQueue.scala 131:72:@10724.4]
  assign _T_10475 = offsetQ_11 < 4'h9; // @[LoadQueue.scala 132:33:@10725.4]
  assign _T_10478 = _T_10475 & _T_6277; // @[LoadQueue.scala 132:41:@10727.4]
  assign _T_10480 = _T_10478 == 1'h0; // @[LoadQueue.scala 132:9:@10728.4]
  assign storesToCheck_11_9 = _T_2558 ? _T_10473 : _T_10480; // @[LoadQueue.scala 131:10:@10729.4]
  assign _T_10486 = 4'ha <= offsetQ_11; // @[LoadQueue.scala 131:81:@10732.4]
  assign _T_10487 = _T_6285 & _T_10486; // @[LoadQueue.scala 131:72:@10733.4]
  assign _T_10489 = offsetQ_11 < 4'ha; // @[LoadQueue.scala 132:33:@10734.4]
  assign _T_10492 = _T_10489 & _T_6294; // @[LoadQueue.scala 132:41:@10736.4]
  assign _T_10494 = _T_10492 == 1'h0; // @[LoadQueue.scala 132:9:@10737.4]
  assign storesToCheck_11_10 = _T_2558 ? _T_10487 : _T_10494; // @[LoadQueue.scala 131:10:@10738.4]
  assign _T_10500 = 4'hb <= offsetQ_11; // @[LoadQueue.scala 131:81:@10741.4]
  assign _T_10501 = _T_6302 & _T_10500; // @[LoadQueue.scala 131:72:@10742.4]
  assign _T_10503 = offsetQ_11 < 4'hb; // @[LoadQueue.scala 132:33:@10743.4]
  assign _T_10506 = _T_10503 & _T_6311; // @[LoadQueue.scala 132:41:@10745.4]
  assign _T_10508 = _T_10506 == 1'h0; // @[LoadQueue.scala 132:9:@10746.4]
  assign storesToCheck_11_11 = _T_2558 ? _T_10501 : _T_10508; // @[LoadQueue.scala 131:10:@10747.4]
  assign _T_10514 = 4'hc <= offsetQ_11; // @[LoadQueue.scala 131:81:@10750.4]
  assign _T_10515 = _T_6319 & _T_10514; // @[LoadQueue.scala 131:72:@10751.4]
  assign _T_10517 = offsetQ_11 < 4'hc; // @[LoadQueue.scala 132:33:@10752.4]
  assign _T_10520 = _T_10517 & _T_6328; // @[LoadQueue.scala 132:41:@10754.4]
  assign _T_10522 = _T_10520 == 1'h0; // @[LoadQueue.scala 132:9:@10755.4]
  assign storesToCheck_11_12 = _T_2558 ? _T_10515 : _T_10522; // @[LoadQueue.scala 131:10:@10756.4]
  assign _T_10528 = 4'hd <= offsetQ_11; // @[LoadQueue.scala 131:81:@10759.4]
  assign _T_10529 = _T_6336 & _T_10528; // @[LoadQueue.scala 131:72:@10760.4]
  assign _T_10531 = offsetQ_11 < 4'hd; // @[LoadQueue.scala 132:33:@10761.4]
  assign _T_10534 = _T_10531 & _T_6345; // @[LoadQueue.scala 132:41:@10763.4]
  assign _T_10536 = _T_10534 == 1'h0; // @[LoadQueue.scala 132:9:@10764.4]
  assign storesToCheck_11_13 = _T_2558 ? _T_10529 : _T_10536; // @[LoadQueue.scala 131:10:@10765.4]
  assign _T_10542 = 4'he <= offsetQ_11; // @[LoadQueue.scala 131:81:@10768.4]
  assign _T_10543 = _T_6353 & _T_10542; // @[LoadQueue.scala 131:72:@10769.4]
  assign _T_10545 = offsetQ_11 < 4'he; // @[LoadQueue.scala 132:33:@10770.4]
  assign _T_10548 = _T_10545 & _T_6362; // @[LoadQueue.scala 132:41:@10772.4]
  assign _T_10550 = _T_10548 == 1'h0; // @[LoadQueue.scala 132:9:@10773.4]
  assign storesToCheck_11_14 = _T_2558 ? _T_10543 : _T_10550; // @[LoadQueue.scala 131:10:@10774.4]
  assign _T_10556 = 4'hf <= offsetQ_11; // @[LoadQueue.scala 131:81:@10777.4]
  assign storesToCheck_11_15 = _T_2558 ? _T_10556 : 1'h1; // @[LoadQueue.scala 131:10:@10783.4]
  assign storesToCheck_12_0 = _T_2588 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@10825.4]
  assign _T_10606 = 4'h1 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10828.4]
  assign _T_10607 = _T_6132 & _T_10606; // @[LoadQueue.scala 131:72:@10829.4]
  assign _T_10609 = offsetQ_12 < 4'h1; // @[LoadQueue.scala 132:33:@10830.4]
  assign _T_10612 = _T_10609 & _T_6141; // @[LoadQueue.scala 132:41:@10832.4]
  assign _T_10614 = _T_10612 == 1'h0; // @[LoadQueue.scala 132:9:@10833.4]
  assign storesToCheck_12_1 = _T_2588 ? _T_10607 : _T_10614; // @[LoadQueue.scala 131:10:@10834.4]
  assign _T_10620 = 4'h2 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10837.4]
  assign _T_10621 = _T_6149 & _T_10620; // @[LoadQueue.scala 131:72:@10838.4]
  assign _T_10623 = offsetQ_12 < 4'h2; // @[LoadQueue.scala 132:33:@10839.4]
  assign _T_10626 = _T_10623 & _T_6158; // @[LoadQueue.scala 132:41:@10841.4]
  assign _T_10628 = _T_10626 == 1'h0; // @[LoadQueue.scala 132:9:@10842.4]
  assign storesToCheck_12_2 = _T_2588 ? _T_10621 : _T_10628; // @[LoadQueue.scala 131:10:@10843.4]
  assign _T_10634 = 4'h3 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10846.4]
  assign _T_10635 = _T_6166 & _T_10634; // @[LoadQueue.scala 131:72:@10847.4]
  assign _T_10637 = offsetQ_12 < 4'h3; // @[LoadQueue.scala 132:33:@10848.4]
  assign _T_10640 = _T_10637 & _T_6175; // @[LoadQueue.scala 132:41:@10850.4]
  assign _T_10642 = _T_10640 == 1'h0; // @[LoadQueue.scala 132:9:@10851.4]
  assign storesToCheck_12_3 = _T_2588 ? _T_10635 : _T_10642; // @[LoadQueue.scala 131:10:@10852.4]
  assign _T_10648 = 4'h4 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10855.4]
  assign _T_10649 = _T_6183 & _T_10648; // @[LoadQueue.scala 131:72:@10856.4]
  assign _T_10651 = offsetQ_12 < 4'h4; // @[LoadQueue.scala 132:33:@10857.4]
  assign _T_10654 = _T_10651 & _T_6192; // @[LoadQueue.scala 132:41:@10859.4]
  assign _T_10656 = _T_10654 == 1'h0; // @[LoadQueue.scala 132:9:@10860.4]
  assign storesToCheck_12_4 = _T_2588 ? _T_10649 : _T_10656; // @[LoadQueue.scala 131:10:@10861.4]
  assign _T_10662 = 4'h5 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10864.4]
  assign _T_10663 = _T_6200 & _T_10662; // @[LoadQueue.scala 131:72:@10865.4]
  assign _T_10665 = offsetQ_12 < 4'h5; // @[LoadQueue.scala 132:33:@10866.4]
  assign _T_10668 = _T_10665 & _T_6209; // @[LoadQueue.scala 132:41:@10868.4]
  assign _T_10670 = _T_10668 == 1'h0; // @[LoadQueue.scala 132:9:@10869.4]
  assign storesToCheck_12_5 = _T_2588 ? _T_10663 : _T_10670; // @[LoadQueue.scala 131:10:@10870.4]
  assign _T_10676 = 4'h6 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10873.4]
  assign _T_10677 = _T_6217 & _T_10676; // @[LoadQueue.scala 131:72:@10874.4]
  assign _T_10679 = offsetQ_12 < 4'h6; // @[LoadQueue.scala 132:33:@10875.4]
  assign _T_10682 = _T_10679 & _T_6226; // @[LoadQueue.scala 132:41:@10877.4]
  assign _T_10684 = _T_10682 == 1'h0; // @[LoadQueue.scala 132:9:@10878.4]
  assign storesToCheck_12_6 = _T_2588 ? _T_10677 : _T_10684; // @[LoadQueue.scala 131:10:@10879.4]
  assign _T_10690 = 4'h7 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10882.4]
  assign _T_10691 = _T_6234 & _T_10690; // @[LoadQueue.scala 131:72:@10883.4]
  assign _T_10693 = offsetQ_12 < 4'h7; // @[LoadQueue.scala 132:33:@10884.4]
  assign _T_10696 = _T_10693 & _T_6243; // @[LoadQueue.scala 132:41:@10886.4]
  assign _T_10698 = _T_10696 == 1'h0; // @[LoadQueue.scala 132:9:@10887.4]
  assign storesToCheck_12_7 = _T_2588 ? _T_10691 : _T_10698; // @[LoadQueue.scala 131:10:@10888.4]
  assign _T_10704 = 4'h8 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10891.4]
  assign _T_10705 = _T_6251 & _T_10704; // @[LoadQueue.scala 131:72:@10892.4]
  assign _T_10707 = offsetQ_12 < 4'h8; // @[LoadQueue.scala 132:33:@10893.4]
  assign _T_10710 = _T_10707 & _T_6260; // @[LoadQueue.scala 132:41:@10895.4]
  assign _T_10712 = _T_10710 == 1'h0; // @[LoadQueue.scala 132:9:@10896.4]
  assign storesToCheck_12_8 = _T_2588 ? _T_10705 : _T_10712; // @[LoadQueue.scala 131:10:@10897.4]
  assign _T_10718 = 4'h9 <= offsetQ_12; // @[LoadQueue.scala 131:81:@10900.4]
  assign _T_10719 = _T_6268 & _T_10718; // @[LoadQueue.scala 131:72:@10901.4]
  assign _T_10721 = offsetQ_12 < 4'h9; // @[LoadQueue.scala 132:33:@10902.4]
  assign _T_10724 = _T_10721 & _T_6277; // @[LoadQueue.scala 132:41:@10904.4]
  assign _T_10726 = _T_10724 == 1'h0; // @[LoadQueue.scala 132:9:@10905.4]
  assign storesToCheck_12_9 = _T_2588 ? _T_10719 : _T_10726; // @[LoadQueue.scala 131:10:@10906.4]
  assign _T_10732 = 4'ha <= offsetQ_12; // @[LoadQueue.scala 131:81:@10909.4]
  assign _T_10733 = _T_6285 & _T_10732; // @[LoadQueue.scala 131:72:@10910.4]
  assign _T_10735 = offsetQ_12 < 4'ha; // @[LoadQueue.scala 132:33:@10911.4]
  assign _T_10738 = _T_10735 & _T_6294; // @[LoadQueue.scala 132:41:@10913.4]
  assign _T_10740 = _T_10738 == 1'h0; // @[LoadQueue.scala 132:9:@10914.4]
  assign storesToCheck_12_10 = _T_2588 ? _T_10733 : _T_10740; // @[LoadQueue.scala 131:10:@10915.4]
  assign _T_10746 = 4'hb <= offsetQ_12; // @[LoadQueue.scala 131:81:@10918.4]
  assign _T_10747 = _T_6302 & _T_10746; // @[LoadQueue.scala 131:72:@10919.4]
  assign _T_10749 = offsetQ_12 < 4'hb; // @[LoadQueue.scala 132:33:@10920.4]
  assign _T_10752 = _T_10749 & _T_6311; // @[LoadQueue.scala 132:41:@10922.4]
  assign _T_10754 = _T_10752 == 1'h0; // @[LoadQueue.scala 132:9:@10923.4]
  assign storesToCheck_12_11 = _T_2588 ? _T_10747 : _T_10754; // @[LoadQueue.scala 131:10:@10924.4]
  assign _T_10760 = 4'hc <= offsetQ_12; // @[LoadQueue.scala 131:81:@10927.4]
  assign _T_10761 = _T_6319 & _T_10760; // @[LoadQueue.scala 131:72:@10928.4]
  assign _T_10763 = offsetQ_12 < 4'hc; // @[LoadQueue.scala 132:33:@10929.4]
  assign _T_10766 = _T_10763 & _T_6328; // @[LoadQueue.scala 132:41:@10931.4]
  assign _T_10768 = _T_10766 == 1'h0; // @[LoadQueue.scala 132:9:@10932.4]
  assign storesToCheck_12_12 = _T_2588 ? _T_10761 : _T_10768; // @[LoadQueue.scala 131:10:@10933.4]
  assign _T_10774 = 4'hd <= offsetQ_12; // @[LoadQueue.scala 131:81:@10936.4]
  assign _T_10775 = _T_6336 & _T_10774; // @[LoadQueue.scala 131:72:@10937.4]
  assign _T_10777 = offsetQ_12 < 4'hd; // @[LoadQueue.scala 132:33:@10938.4]
  assign _T_10780 = _T_10777 & _T_6345; // @[LoadQueue.scala 132:41:@10940.4]
  assign _T_10782 = _T_10780 == 1'h0; // @[LoadQueue.scala 132:9:@10941.4]
  assign storesToCheck_12_13 = _T_2588 ? _T_10775 : _T_10782; // @[LoadQueue.scala 131:10:@10942.4]
  assign _T_10788 = 4'he <= offsetQ_12; // @[LoadQueue.scala 131:81:@10945.4]
  assign _T_10789 = _T_6353 & _T_10788; // @[LoadQueue.scala 131:72:@10946.4]
  assign _T_10791 = offsetQ_12 < 4'he; // @[LoadQueue.scala 132:33:@10947.4]
  assign _T_10794 = _T_10791 & _T_6362; // @[LoadQueue.scala 132:41:@10949.4]
  assign _T_10796 = _T_10794 == 1'h0; // @[LoadQueue.scala 132:9:@10950.4]
  assign storesToCheck_12_14 = _T_2588 ? _T_10789 : _T_10796; // @[LoadQueue.scala 131:10:@10951.4]
  assign _T_10802 = 4'hf <= offsetQ_12; // @[LoadQueue.scala 131:81:@10954.4]
  assign storesToCheck_12_15 = _T_2588 ? _T_10802 : 1'h1; // @[LoadQueue.scala 131:10:@10960.4]
  assign storesToCheck_13_0 = _T_2618 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11002.4]
  assign _T_10852 = 4'h1 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11005.4]
  assign _T_10853 = _T_6132 & _T_10852; // @[LoadQueue.scala 131:72:@11006.4]
  assign _T_10855 = offsetQ_13 < 4'h1; // @[LoadQueue.scala 132:33:@11007.4]
  assign _T_10858 = _T_10855 & _T_6141; // @[LoadQueue.scala 132:41:@11009.4]
  assign _T_10860 = _T_10858 == 1'h0; // @[LoadQueue.scala 132:9:@11010.4]
  assign storesToCheck_13_1 = _T_2618 ? _T_10853 : _T_10860; // @[LoadQueue.scala 131:10:@11011.4]
  assign _T_10866 = 4'h2 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11014.4]
  assign _T_10867 = _T_6149 & _T_10866; // @[LoadQueue.scala 131:72:@11015.4]
  assign _T_10869 = offsetQ_13 < 4'h2; // @[LoadQueue.scala 132:33:@11016.4]
  assign _T_10872 = _T_10869 & _T_6158; // @[LoadQueue.scala 132:41:@11018.4]
  assign _T_10874 = _T_10872 == 1'h0; // @[LoadQueue.scala 132:9:@11019.4]
  assign storesToCheck_13_2 = _T_2618 ? _T_10867 : _T_10874; // @[LoadQueue.scala 131:10:@11020.4]
  assign _T_10880 = 4'h3 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11023.4]
  assign _T_10881 = _T_6166 & _T_10880; // @[LoadQueue.scala 131:72:@11024.4]
  assign _T_10883 = offsetQ_13 < 4'h3; // @[LoadQueue.scala 132:33:@11025.4]
  assign _T_10886 = _T_10883 & _T_6175; // @[LoadQueue.scala 132:41:@11027.4]
  assign _T_10888 = _T_10886 == 1'h0; // @[LoadQueue.scala 132:9:@11028.4]
  assign storesToCheck_13_3 = _T_2618 ? _T_10881 : _T_10888; // @[LoadQueue.scala 131:10:@11029.4]
  assign _T_10894 = 4'h4 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11032.4]
  assign _T_10895 = _T_6183 & _T_10894; // @[LoadQueue.scala 131:72:@11033.4]
  assign _T_10897 = offsetQ_13 < 4'h4; // @[LoadQueue.scala 132:33:@11034.4]
  assign _T_10900 = _T_10897 & _T_6192; // @[LoadQueue.scala 132:41:@11036.4]
  assign _T_10902 = _T_10900 == 1'h0; // @[LoadQueue.scala 132:9:@11037.4]
  assign storesToCheck_13_4 = _T_2618 ? _T_10895 : _T_10902; // @[LoadQueue.scala 131:10:@11038.4]
  assign _T_10908 = 4'h5 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11041.4]
  assign _T_10909 = _T_6200 & _T_10908; // @[LoadQueue.scala 131:72:@11042.4]
  assign _T_10911 = offsetQ_13 < 4'h5; // @[LoadQueue.scala 132:33:@11043.4]
  assign _T_10914 = _T_10911 & _T_6209; // @[LoadQueue.scala 132:41:@11045.4]
  assign _T_10916 = _T_10914 == 1'h0; // @[LoadQueue.scala 132:9:@11046.4]
  assign storesToCheck_13_5 = _T_2618 ? _T_10909 : _T_10916; // @[LoadQueue.scala 131:10:@11047.4]
  assign _T_10922 = 4'h6 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11050.4]
  assign _T_10923 = _T_6217 & _T_10922; // @[LoadQueue.scala 131:72:@11051.4]
  assign _T_10925 = offsetQ_13 < 4'h6; // @[LoadQueue.scala 132:33:@11052.4]
  assign _T_10928 = _T_10925 & _T_6226; // @[LoadQueue.scala 132:41:@11054.4]
  assign _T_10930 = _T_10928 == 1'h0; // @[LoadQueue.scala 132:9:@11055.4]
  assign storesToCheck_13_6 = _T_2618 ? _T_10923 : _T_10930; // @[LoadQueue.scala 131:10:@11056.4]
  assign _T_10936 = 4'h7 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11059.4]
  assign _T_10937 = _T_6234 & _T_10936; // @[LoadQueue.scala 131:72:@11060.4]
  assign _T_10939 = offsetQ_13 < 4'h7; // @[LoadQueue.scala 132:33:@11061.4]
  assign _T_10942 = _T_10939 & _T_6243; // @[LoadQueue.scala 132:41:@11063.4]
  assign _T_10944 = _T_10942 == 1'h0; // @[LoadQueue.scala 132:9:@11064.4]
  assign storesToCheck_13_7 = _T_2618 ? _T_10937 : _T_10944; // @[LoadQueue.scala 131:10:@11065.4]
  assign _T_10950 = 4'h8 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11068.4]
  assign _T_10951 = _T_6251 & _T_10950; // @[LoadQueue.scala 131:72:@11069.4]
  assign _T_10953 = offsetQ_13 < 4'h8; // @[LoadQueue.scala 132:33:@11070.4]
  assign _T_10956 = _T_10953 & _T_6260; // @[LoadQueue.scala 132:41:@11072.4]
  assign _T_10958 = _T_10956 == 1'h0; // @[LoadQueue.scala 132:9:@11073.4]
  assign storesToCheck_13_8 = _T_2618 ? _T_10951 : _T_10958; // @[LoadQueue.scala 131:10:@11074.4]
  assign _T_10964 = 4'h9 <= offsetQ_13; // @[LoadQueue.scala 131:81:@11077.4]
  assign _T_10965 = _T_6268 & _T_10964; // @[LoadQueue.scala 131:72:@11078.4]
  assign _T_10967 = offsetQ_13 < 4'h9; // @[LoadQueue.scala 132:33:@11079.4]
  assign _T_10970 = _T_10967 & _T_6277; // @[LoadQueue.scala 132:41:@11081.4]
  assign _T_10972 = _T_10970 == 1'h0; // @[LoadQueue.scala 132:9:@11082.4]
  assign storesToCheck_13_9 = _T_2618 ? _T_10965 : _T_10972; // @[LoadQueue.scala 131:10:@11083.4]
  assign _T_10978 = 4'ha <= offsetQ_13; // @[LoadQueue.scala 131:81:@11086.4]
  assign _T_10979 = _T_6285 & _T_10978; // @[LoadQueue.scala 131:72:@11087.4]
  assign _T_10981 = offsetQ_13 < 4'ha; // @[LoadQueue.scala 132:33:@11088.4]
  assign _T_10984 = _T_10981 & _T_6294; // @[LoadQueue.scala 132:41:@11090.4]
  assign _T_10986 = _T_10984 == 1'h0; // @[LoadQueue.scala 132:9:@11091.4]
  assign storesToCheck_13_10 = _T_2618 ? _T_10979 : _T_10986; // @[LoadQueue.scala 131:10:@11092.4]
  assign _T_10992 = 4'hb <= offsetQ_13; // @[LoadQueue.scala 131:81:@11095.4]
  assign _T_10993 = _T_6302 & _T_10992; // @[LoadQueue.scala 131:72:@11096.4]
  assign _T_10995 = offsetQ_13 < 4'hb; // @[LoadQueue.scala 132:33:@11097.4]
  assign _T_10998 = _T_10995 & _T_6311; // @[LoadQueue.scala 132:41:@11099.4]
  assign _T_11000 = _T_10998 == 1'h0; // @[LoadQueue.scala 132:9:@11100.4]
  assign storesToCheck_13_11 = _T_2618 ? _T_10993 : _T_11000; // @[LoadQueue.scala 131:10:@11101.4]
  assign _T_11006 = 4'hc <= offsetQ_13; // @[LoadQueue.scala 131:81:@11104.4]
  assign _T_11007 = _T_6319 & _T_11006; // @[LoadQueue.scala 131:72:@11105.4]
  assign _T_11009 = offsetQ_13 < 4'hc; // @[LoadQueue.scala 132:33:@11106.4]
  assign _T_11012 = _T_11009 & _T_6328; // @[LoadQueue.scala 132:41:@11108.4]
  assign _T_11014 = _T_11012 == 1'h0; // @[LoadQueue.scala 132:9:@11109.4]
  assign storesToCheck_13_12 = _T_2618 ? _T_11007 : _T_11014; // @[LoadQueue.scala 131:10:@11110.4]
  assign _T_11020 = 4'hd <= offsetQ_13; // @[LoadQueue.scala 131:81:@11113.4]
  assign _T_11021 = _T_6336 & _T_11020; // @[LoadQueue.scala 131:72:@11114.4]
  assign _T_11023 = offsetQ_13 < 4'hd; // @[LoadQueue.scala 132:33:@11115.4]
  assign _T_11026 = _T_11023 & _T_6345; // @[LoadQueue.scala 132:41:@11117.4]
  assign _T_11028 = _T_11026 == 1'h0; // @[LoadQueue.scala 132:9:@11118.4]
  assign storesToCheck_13_13 = _T_2618 ? _T_11021 : _T_11028; // @[LoadQueue.scala 131:10:@11119.4]
  assign _T_11034 = 4'he <= offsetQ_13; // @[LoadQueue.scala 131:81:@11122.4]
  assign _T_11035 = _T_6353 & _T_11034; // @[LoadQueue.scala 131:72:@11123.4]
  assign _T_11037 = offsetQ_13 < 4'he; // @[LoadQueue.scala 132:33:@11124.4]
  assign _T_11040 = _T_11037 & _T_6362; // @[LoadQueue.scala 132:41:@11126.4]
  assign _T_11042 = _T_11040 == 1'h0; // @[LoadQueue.scala 132:9:@11127.4]
  assign storesToCheck_13_14 = _T_2618 ? _T_11035 : _T_11042; // @[LoadQueue.scala 131:10:@11128.4]
  assign _T_11048 = 4'hf <= offsetQ_13; // @[LoadQueue.scala 131:81:@11131.4]
  assign storesToCheck_13_15 = _T_2618 ? _T_11048 : 1'h1; // @[LoadQueue.scala 131:10:@11137.4]
  assign storesToCheck_14_0 = _T_2648 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11179.4]
  assign _T_11098 = 4'h1 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11182.4]
  assign _T_11099 = _T_6132 & _T_11098; // @[LoadQueue.scala 131:72:@11183.4]
  assign _T_11101 = offsetQ_14 < 4'h1; // @[LoadQueue.scala 132:33:@11184.4]
  assign _T_11104 = _T_11101 & _T_6141; // @[LoadQueue.scala 132:41:@11186.4]
  assign _T_11106 = _T_11104 == 1'h0; // @[LoadQueue.scala 132:9:@11187.4]
  assign storesToCheck_14_1 = _T_2648 ? _T_11099 : _T_11106; // @[LoadQueue.scala 131:10:@11188.4]
  assign _T_11112 = 4'h2 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11191.4]
  assign _T_11113 = _T_6149 & _T_11112; // @[LoadQueue.scala 131:72:@11192.4]
  assign _T_11115 = offsetQ_14 < 4'h2; // @[LoadQueue.scala 132:33:@11193.4]
  assign _T_11118 = _T_11115 & _T_6158; // @[LoadQueue.scala 132:41:@11195.4]
  assign _T_11120 = _T_11118 == 1'h0; // @[LoadQueue.scala 132:9:@11196.4]
  assign storesToCheck_14_2 = _T_2648 ? _T_11113 : _T_11120; // @[LoadQueue.scala 131:10:@11197.4]
  assign _T_11126 = 4'h3 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11200.4]
  assign _T_11127 = _T_6166 & _T_11126; // @[LoadQueue.scala 131:72:@11201.4]
  assign _T_11129 = offsetQ_14 < 4'h3; // @[LoadQueue.scala 132:33:@11202.4]
  assign _T_11132 = _T_11129 & _T_6175; // @[LoadQueue.scala 132:41:@11204.4]
  assign _T_11134 = _T_11132 == 1'h0; // @[LoadQueue.scala 132:9:@11205.4]
  assign storesToCheck_14_3 = _T_2648 ? _T_11127 : _T_11134; // @[LoadQueue.scala 131:10:@11206.4]
  assign _T_11140 = 4'h4 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11209.4]
  assign _T_11141 = _T_6183 & _T_11140; // @[LoadQueue.scala 131:72:@11210.4]
  assign _T_11143 = offsetQ_14 < 4'h4; // @[LoadQueue.scala 132:33:@11211.4]
  assign _T_11146 = _T_11143 & _T_6192; // @[LoadQueue.scala 132:41:@11213.4]
  assign _T_11148 = _T_11146 == 1'h0; // @[LoadQueue.scala 132:9:@11214.4]
  assign storesToCheck_14_4 = _T_2648 ? _T_11141 : _T_11148; // @[LoadQueue.scala 131:10:@11215.4]
  assign _T_11154 = 4'h5 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11218.4]
  assign _T_11155 = _T_6200 & _T_11154; // @[LoadQueue.scala 131:72:@11219.4]
  assign _T_11157 = offsetQ_14 < 4'h5; // @[LoadQueue.scala 132:33:@11220.4]
  assign _T_11160 = _T_11157 & _T_6209; // @[LoadQueue.scala 132:41:@11222.4]
  assign _T_11162 = _T_11160 == 1'h0; // @[LoadQueue.scala 132:9:@11223.4]
  assign storesToCheck_14_5 = _T_2648 ? _T_11155 : _T_11162; // @[LoadQueue.scala 131:10:@11224.4]
  assign _T_11168 = 4'h6 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11227.4]
  assign _T_11169 = _T_6217 & _T_11168; // @[LoadQueue.scala 131:72:@11228.4]
  assign _T_11171 = offsetQ_14 < 4'h6; // @[LoadQueue.scala 132:33:@11229.4]
  assign _T_11174 = _T_11171 & _T_6226; // @[LoadQueue.scala 132:41:@11231.4]
  assign _T_11176 = _T_11174 == 1'h0; // @[LoadQueue.scala 132:9:@11232.4]
  assign storesToCheck_14_6 = _T_2648 ? _T_11169 : _T_11176; // @[LoadQueue.scala 131:10:@11233.4]
  assign _T_11182 = 4'h7 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11236.4]
  assign _T_11183 = _T_6234 & _T_11182; // @[LoadQueue.scala 131:72:@11237.4]
  assign _T_11185 = offsetQ_14 < 4'h7; // @[LoadQueue.scala 132:33:@11238.4]
  assign _T_11188 = _T_11185 & _T_6243; // @[LoadQueue.scala 132:41:@11240.4]
  assign _T_11190 = _T_11188 == 1'h0; // @[LoadQueue.scala 132:9:@11241.4]
  assign storesToCheck_14_7 = _T_2648 ? _T_11183 : _T_11190; // @[LoadQueue.scala 131:10:@11242.4]
  assign _T_11196 = 4'h8 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11245.4]
  assign _T_11197 = _T_6251 & _T_11196; // @[LoadQueue.scala 131:72:@11246.4]
  assign _T_11199 = offsetQ_14 < 4'h8; // @[LoadQueue.scala 132:33:@11247.4]
  assign _T_11202 = _T_11199 & _T_6260; // @[LoadQueue.scala 132:41:@11249.4]
  assign _T_11204 = _T_11202 == 1'h0; // @[LoadQueue.scala 132:9:@11250.4]
  assign storesToCheck_14_8 = _T_2648 ? _T_11197 : _T_11204; // @[LoadQueue.scala 131:10:@11251.4]
  assign _T_11210 = 4'h9 <= offsetQ_14; // @[LoadQueue.scala 131:81:@11254.4]
  assign _T_11211 = _T_6268 & _T_11210; // @[LoadQueue.scala 131:72:@11255.4]
  assign _T_11213 = offsetQ_14 < 4'h9; // @[LoadQueue.scala 132:33:@11256.4]
  assign _T_11216 = _T_11213 & _T_6277; // @[LoadQueue.scala 132:41:@11258.4]
  assign _T_11218 = _T_11216 == 1'h0; // @[LoadQueue.scala 132:9:@11259.4]
  assign storesToCheck_14_9 = _T_2648 ? _T_11211 : _T_11218; // @[LoadQueue.scala 131:10:@11260.4]
  assign _T_11224 = 4'ha <= offsetQ_14; // @[LoadQueue.scala 131:81:@11263.4]
  assign _T_11225 = _T_6285 & _T_11224; // @[LoadQueue.scala 131:72:@11264.4]
  assign _T_11227 = offsetQ_14 < 4'ha; // @[LoadQueue.scala 132:33:@11265.4]
  assign _T_11230 = _T_11227 & _T_6294; // @[LoadQueue.scala 132:41:@11267.4]
  assign _T_11232 = _T_11230 == 1'h0; // @[LoadQueue.scala 132:9:@11268.4]
  assign storesToCheck_14_10 = _T_2648 ? _T_11225 : _T_11232; // @[LoadQueue.scala 131:10:@11269.4]
  assign _T_11238 = 4'hb <= offsetQ_14; // @[LoadQueue.scala 131:81:@11272.4]
  assign _T_11239 = _T_6302 & _T_11238; // @[LoadQueue.scala 131:72:@11273.4]
  assign _T_11241 = offsetQ_14 < 4'hb; // @[LoadQueue.scala 132:33:@11274.4]
  assign _T_11244 = _T_11241 & _T_6311; // @[LoadQueue.scala 132:41:@11276.4]
  assign _T_11246 = _T_11244 == 1'h0; // @[LoadQueue.scala 132:9:@11277.4]
  assign storesToCheck_14_11 = _T_2648 ? _T_11239 : _T_11246; // @[LoadQueue.scala 131:10:@11278.4]
  assign _T_11252 = 4'hc <= offsetQ_14; // @[LoadQueue.scala 131:81:@11281.4]
  assign _T_11253 = _T_6319 & _T_11252; // @[LoadQueue.scala 131:72:@11282.4]
  assign _T_11255 = offsetQ_14 < 4'hc; // @[LoadQueue.scala 132:33:@11283.4]
  assign _T_11258 = _T_11255 & _T_6328; // @[LoadQueue.scala 132:41:@11285.4]
  assign _T_11260 = _T_11258 == 1'h0; // @[LoadQueue.scala 132:9:@11286.4]
  assign storesToCheck_14_12 = _T_2648 ? _T_11253 : _T_11260; // @[LoadQueue.scala 131:10:@11287.4]
  assign _T_11266 = 4'hd <= offsetQ_14; // @[LoadQueue.scala 131:81:@11290.4]
  assign _T_11267 = _T_6336 & _T_11266; // @[LoadQueue.scala 131:72:@11291.4]
  assign _T_11269 = offsetQ_14 < 4'hd; // @[LoadQueue.scala 132:33:@11292.4]
  assign _T_11272 = _T_11269 & _T_6345; // @[LoadQueue.scala 132:41:@11294.4]
  assign _T_11274 = _T_11272 == 1'h0; // @[LoadQueue.scala 132:9:@11295.4]
  assign storesToCheck_14_13 = _T_2648 ? _T_11267 : _T_11274; // @[LoadQueue.scala 131:10:@11296.4]
  assign _T_11280 = 4'he <= offsetQ_14; // @[LoadQueue.scala 131:81:@11299.4]
  assign _T_11281 = _T_6353 & _T_11280; // @[LoadQueue.scala 131:72:@11300.4]
  assign _T_11283 = offsetQ_14 < 4'he; // @[LoadQueue.scala 132:33:@11301.4]
  assign _T_11286 = _T_11283 & _T_6362; // @[LoadQueue.scala 132:41:@11303.4]
  assign _T_11288 = _T_11286 == 1'h0; // @[LoadQueue.scala 132:9:@11304.4]
  assign storesToCheck_14_14 = _T_2648 ? _T_11281 : _T_11288; // @[LoadQueue.scala 131:10:@11305.4]
  assign _T_11294 = 4'hf <= offsetQ_14; // @[LoadQueue.scala 131:81:@11308.4]
  assign storesToCheck_14_15 = _T_2648 ? _T_11294 : 1'h1; // @[LoadQueue.scala 131:10:@11314.4]
  assign storesToCheck_15_0 = _T_2678 ? _T_6115 : 1'h1; // @[LoadQueue.scala 131:10:@11356.4]
  assign _T_11344 = 4'h1 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11359.4]
  assign _T_11345 = _T_6132 & _T_11344; // @[LoadQueue.scala 131:72:@11360.4]
  assign _T_11347 = offsetQ_15 < 4'h1; // @[LoadQueue.scala 132:33:@11361.4]
  assign _T_11350 = _T_11347 & _T_6141; // @[LoadQueue.scala 132:41:@11363.4]
  assign _T_11352 = _T_11350 == 1'h0; // @[LoadQueue.scala 132:9:@11364.4]
  assign storesToCheck_15_1 = _T_2678 ? _T_11345 : _T_11352; // @[LoadQueue.scala 131:10:@11365.4]
  assign _T_11358 = 4'h2 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11368.4]
  assign _T_11359 = _T_6149 & _T_11358; // @[LoadQueue.scala 131:72:@11369.4]
  assign _T_11361 = offsetQ_15 < 4'h2; // @[LoadQueue.scala 132:33:@11370.4]
  assign _T_11364 = _T_11361 & _T_6158; // @[LoadQueue.scala 132:41:@11372.4]
  assign _T_11366 = _T_11364 == 1'h0; // @[LoadQueue.scala 132:9:@11373.4]
  assign storesToCheck_15_2 = _T_2678 ? _T_11359 : _T_11366; // @[LoadQueue.scala 131:10:@11374.4]
  assign _T_11372 = 4'h3 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11377.4]
  assign _T_11373 = _T_6166 & _T_11372; // @[LoadQueue.scala 131:72:@11378.4]
  assign _T_11375 = offsetQ_15 < 4'h3; // @[LoadQueue.scala 132:33:@11379.4]
  assign _T_11378 = _T_11375 & _T_6175; // @[LoadQueue.scala 132:41:@11381.4]
  assign _T_11380 = _T_11378 == 1'h0; // @[LoadQueue.scala 132:9:@11382.4]
  assign storesToCheck_15_3 = _T_2678 ? _T_11373 : _T_11380; // @[LoadQueue.scala 131:10:@11383.4]
  assign _T_11386 = 4'h4 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11386.4]
  assign _T_11387 = _T_6183 & _T_11386; // @[LoadQueue.scala 131:72:@11387.4]
  assign _T_11389 = offsetQ_15 < 4'h4; // @[LoadQueue.scala 132:33:@11388.4]
  assign _T_11392 = _T_11389 & _T_6192; // @[LoadQueue.scala 132:41:@11390.4]
  assign _T_11394 = _T_11392 == 1'h0; // @[LoadQueue.scala 132:9:@11391.4]
  assign storesToCheck_15_4 = _T_2678 ? _T_11387 : _T_11394; // @[LoadQueue.scala 131:10:@11392.4]
  assign _T_11400 = 4'h5 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11395.4]
  assign _T_11401 = _T_6200 & _T_11400; // @[LoadQueue.scala 131:72:@11396.4]
  assign _T_11403 = offsetQ_15 < 4'h5; // @[LoadQueue.scala 132:33:@11397.4]
  assign _T_11406 = _T_11403 & _T_6209; // @[LoadQueue.scala 132:41:@11399.4]
  assign _T_11408 = _T_11406 == 1'h0; // @[LoadQueue.scala 132:9:@11400.4]
  assign storesToCheck_15_5 = _T_2678 ? _T_11401 : _T_11408; // @[LoadQueue.scala 131:10:@11401.4]
  assign _T_11414 = 4'h6 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11404.4]
  assign _T_11415 = _T_6217 & _T_11414; // @[LoadQueue.scala 131:72:@11405.4]
  assign _T_11417 = offsetQ_15 < 4'h6; // @[LoadQueue.scala 132:33:@11406.4]
  assign _T_11420 = _T_11417 & _T_6226; // @[LoadQueue.scala 132:41:@11408.4]
  assign _T_11422 = _T_11420 == 1'h0; // @[LoadQueue.scala 132:9:@11409.4]
  assign storesToCheck_15_6 = _T_2678 ? _T_11415 : _T_11422; // @[LoadQueue.scala 131:10:@11410.4]
  assign _T_11428 = 4'h7 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11413.4]
  assign _T_11429 = _T_6234 & _T_11428; // @[LoadQueue.scala 131:72:@11414.4]
  assign _T_11431 = offsetQ_15 < 4'h7; // @[LoadQueue.scala 132:33:@11415.4]
  assign _T_11434 = _T_11431 & _T_6243; // @[LoadQueue.scala 132:41:@11417.4]
  assign _T_11436 = _T_11434 == 1'h0; // @[LoadQueue.scala 132:9:@11418.4]
  assign storesToCheck_15_7 = _T_2678 ? _T_11429 : _T_11436; // @[LoadQueue.scala 131:10:@11419.4]
  assign _T_11442 = 4'h8 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11422.4]
  assign _T_11443 = _T_6251 & _T_11442; // @[LoadQueue.scala 131:72:@11423.4]
  assign _T_11445 = offsetQ_15 < 4'h8; // @[LoadQueue.scala 132:33:@11424.4]
  assign _T_11448 = _T_11445 & _T_6260; // @[LoadQueue.scala 132:41:@11426.4]
  assign _T_11450 = _T_11448 == 1'h0; // @[LoadQueue.scala 132:9:@11427.4]
  assign storesToCheck_15_8 = _T_2678 ? _T_11443 : _T_11450; // @[LoadQueue.scala 131:10:@11428.4]
  assign _T_11456 = 4'h9 <= offsetQ_15; // @[LoadQueue.scala 131:81:@11431.4]
  assign _T_11457 = _T_6268 & _T_11456; // @[LoadQueue.scala 131:72:@11432.4]
  assign _T_11459 = offsetQ_15 < 4'h9; // @[LoadQueue.scala 132:33:@11433.4]
  assign _T_11462 = _T_11459 & _T_6277; // @[LoadQueue.scala 132:41:@11435.4]
  assign _T_11464 = _T_11462 == 1'h0; // @[LoadQueue.scala 132:9:@11436.4]
  assign storesToCheck_15_9 = _T_2678 ? _T_11457 : _T_11464; // @[LoadQueue.scala 131:10:@11437.4]
  assign _T_11470 = 4'ha <= offsetQ_15; // @[LoadQueue.scala 131:81:@11440.4]
  assign _T_11471 = _T_6285 & _T_11470; // @[LoadQueue.scala 131:72:@11441.4]
  assign _T_11473 = offsetQ_15 < 4'ha; // @[LoadQueue.scala 132:33:@11442.4]
  assign _T_11476 = _T_11473 & _T_6294; // @[LoadQueue.scala 132:41:@11444.4]
  assign _T_11478 = _T_11476 == 1'h0; // @[LoadQueue.scala 132:9:@11445.4]
  assign storesToCheck_15_10 = _T_2678 ? _T_11471 : _T_11478; // @[LoadQueue.scala 131:10:@11446.4]
  assign _T_11484 = 4'hb <= offsetQ_15; // @[LoadQueue.scala 131:81:@11449.4]
  assign _T_11485 = _T_6302 & _T_11484; // @[LoadQueue.scala 131:72:@11450.4]
  assign _T_11487 = offsetQ_15 < 4'hb; // @[LoadQueue.scala 132:33:@11451.4]
  assign _T_11490 = _T_11487 & _T_6311; // @[LoadQueue.scala 132:41:@11453.4]
  assign _T_11492 = _T_11490 == 1'h0; // @[LoadQueue.scala 132:9:@11454.4]
  assign storesToCheck_15_11 = _T_2678 ? _T_11485 : _T_11492; // @[LoadQueue.scala 131:10:@11455.4]
  assign _T_11498 = 4'hc <= offsetQ_15; // @[LoadQueue.scala 131:81:@11458.4]
  assign _T_11499 = _T_6319 & _T_11498; // @[LoadQueue.scala 131:72:@11459.4]
  assign _T_11501 = offsetQ_15 < 4'hc; // @[LoadQueue.scala 132:33:@11460.4]
  assign _T_11504 = _T_11501 & _T_6328; // @[LoadQueue.scala 132:41:@11462.4]
  assign _T_11506 = _T_11504 == 1'h0; // @[LoadQueue.scala 132:9:@11463.4]
  assign storesToCheck_15_12 = _T_2678 ? _T_11499 : _T_11506; // @[LoadQueue.scala 131:10:@11464.4]
  assign _T_11512 = 4'hd <= offsetQ_15; // @[LoadQueue.scala 131:81:@11467.4]
  assign _T_11513 = _T_6336 & _T_11512; // @[LoadQueue.scala 131:72:@11468.4]
  assign _T_11515 = offsetQ_15 < 4'hd; // @[LoadQueue.scala 132:33:@11469.4]
  assign _T_11518 = _T_11515 & _T_6345; // @[LoadQueue.scala 132:41:@11471.4]
  assign _T_11520 = _T_11518 == 1'h0; // @[LoadQueue.scala 132:9:@11472.4]
  assign storesToCheck_15_13 = _T_2678 ? _T_11513 : _T_11520; // @[LoadQueue.scala 131:10:@11473.4]
  assign _T_11526 = 4'he <= offsetQ_15; // @[LoadQueue.scala 131:81:@11476.4]
  assign _T_11527 = _T_6353 & _T_11526; // @[LoadQueue.scala 131:72:@11477.4]
  assign _T_11529 = offsetQ_15 < 4'he; // @[LoadQueue.scala 132:33:@11478.4]
  assign _T_11532 = _T_11529 & _T_6362; // @[LoadQueue.scala 132:41:@11480.4]
  assign _T_11534 = _T_11532 == 1'h0; // @[LoadQueue.scala 132:9:@11481.4]
  assign storesToCheck_15_14 = _T_2678 ? _T_11527 : _T_11534; // @[LoadQueue.scala 131:10:@11482.4]
  assign _T_11540 = 4'hf <= offsetQ_15; // @[LoadQueue.scala 131:81:@11485.4]
  assign storesToCheck_15_15 = _T_2678 ? _T_11540 : 1'h1; // @[LoadQueue.scala 131:10:@11491.4]
  assign _T_12802 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11526.4]
  assign entriesToCheck_0_0 = _T_12802 & checkBits_0; // @[LoadQueue.scala 141:26:@11527.4]
  assign _T_12804 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11528.4]
  assign entriesToCheck_0_1 = _T_12804 & checkBits_0; // @[LoadQueue.scala 141:26:@11529.4]
  assign _T_12806 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11530.4]
  assign entriesToCheck_0_2 = _T_12806 & checkBits_0; // @[LoadQueue.scala 141:26:@11531.4]
  assign _T_12808 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11532.4]
  assign entriesToCheck_0_3 = _T_12808 & checkBits_0; // @[LoadQueue.scala 141:26:@11533.4]
  assign _T_12810 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11534.4]
  assign entriesToCheck_0_4 = _T_12810 & checkBits_0; // @[LoadQueue.scala 141:26:@11535.4]
  assign _T_12812 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11536.4]
  assign entriesToCheck_0_5 = _T_12812 & checkBits_0; // @[LoadQueue.scala 141:26:@11537.4]
  assign _T_12814 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11538.4]
  assign entriesToCheck_0_6 = _T_12814 & checkBits_0; // @[LoadQueue.scala 141:26:@11539.4]
  assign _T_12816 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11540.4]
  assign entriesToCheck_0_7 = _T_12816 & checkBits_0; // @[LoadQueue.scala 141:26:@11541.4]
  assign _T_12818 = storesToCheck_0_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11542.4]
  assign entriesToCheck_0_8 = _T_12818 & checkBits_0; // @[LoadQueue.scala 141:26:@11543.4]
  assign _T_12820 = storesToCheck_0_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11544.4]
  assign entriesToCheck_0_9 = _T_12820 & checkBits_0; // @[LoadQueue.scala 141:26:@11545.4]
  assign _T_12822 = storesToCheck_0_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11546.4]
  assign entriesToCheck_0_10 = _T_12822 & checkBits_0; // @[LoadQueue.scala 141:26:@11547.4]
  assign _T_12824 = storesToCheck_0_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11548.4]
  assign entriesToCheck_0_11 = _T_12824 & checkBits_0; // @[LoadQueue.scala 141:26:@11549.4]
  assign _T_12826 = storesToCheck_0_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11550.4]
  assign entriesToCheck_0_12 = _T_12826 & checkBits_0; // @[LoadQueue.scala 141:26:@11551.4]
  assign _T_12828 = storesToCheck_0_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11552.4]
  assign entriesToCheck_0_13 = _T_12828 & checkBits_0; // @[LoadQueue.scala 141:26:@11553.4]
  assign _T_12830 = storesToCheck_0_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11554.4]
  assign entriesToCheck_0_14 = _T_12830 & checkBits_0; // @[LoadQueue.scala 141:26:@11555.4]
  assign _T_12832 = storesToCheck_0_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11556.4]
  assign entriesToCheck_0_15 = _T_12832 & checkBits_0; // @[LoadQueue.scala 141:26:@11557.4]
  assign _T_12834 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11574.4]
  assign entriesToCheck_1_0 = _T_12834 & checkBits_1; // @[LoadQueue.scala 141:26:@11575.4]
  assign _T_12836 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11576.4]
  assign entriesToCheck_1_1 = _T_12836 & checkBits_1; // @[LoadQueue.scala 141:26:@11577.4]
  assign _T_12838 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11578.4]
  assign entriesToCheck_1_2 = _T_12838 & checkBits_1; // @[LoadQueue.scala 141:26:@11579.4]
  assign _T_12840 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11580.4]
  assign entriesToCheck_1_3 = _T_12840 & checkBits_1; // @[LoadQueue.scala 141:26:@11581.4]
  assign _T_12842 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11582.4]
  assign entriesToCheck_1_4 = _T_12842 & checkBits_1; // @[LoadQueue.scala 141:26:@11583.4]
  assign _T_12844 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11584.4]
  assign entriesToCheck_1_5 = _T_12844 & checkBits_1; // @[LoadQueue.scala 141:26:@11585.4]
  assign _T_12846 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11586.4]
  assign entriesToCheck_1_6 = _T_12846 & checkBits_1; // @[LoadQueue.scala 141:26:@11587.4]
  assign _T_12848 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11588.4]
  assign entriesToCheck_1_7 = _T_12848 & checkBits_1; // @[LoadQueue.scala 141:26:@11589.4]
  assign _T_12850 = storesToCheck_1_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11590.4]
  assign entriesToCheck_1_8 = _T_12850 & checkBits_1; // @[LoadQueue.scala 141:26:@11591.4]
  assign _T_12852 = storesToCheck_1_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11592.4]
  assign entriesToCheck_1_9 = _T_12852 & checkBits_1; // @[LoadQueue.scala 141:26:@11593.4]
  assign _T_12854 = storesToCheck_1_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11594.4]
  assign entriesToCheck_1_10 = _T_12854 & checkBits_1; // @[LoadQueue.scala 141:26:@11595.4]
  assign _T_12856 = storesToCheck_1_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11596.4]
  assign entriesToCheck_1_11 = _T_12856 & checkBits_1; // @[LoadQueue.scala 141:26:@11597.4]
  assign _T_12858 = storesToCheck_1_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11598.4]
  assign entriesToCheck_1_12 = _T_12858 & checkBits_1; // @[LoadQueue.scala 141:26:@11599.4]
  assign _T_12860 = storesToCheck_1_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11600.4]
  assign entriesToCheck_1_13 = _T_12860 & checkBits_1; // @[LoadQueue.scala 141:26:@11601.4]
  assign _T_12862 = storesToCheck_1_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11602.4]
  assign entriesToCheck_1_14 = _T_12862 & checkBits_1; // @[LoadQueue.scala 141:26:@11603.4]
  assign _T_12864 = storesToCheck_1_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11604.4]
  assign entriesToCheck_1_15 = _T_12864 & checkBits_1; // @[LoadQueue.scala 141:26:@11605.4]
  assign _T_12866 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11622.4]
  assign entriesToCheck_2_0 = _T_12866 & checkBits_2; // @[LoadQueue.scala 141:26:@11623.4]
  assign _T_12868 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11624.4]
  assign entriesToCheck_2_1 = _T_12868 & checkBits_2; // @[LoadQueue.scala 141:26:@11625.4]
  assign _T_12870 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11626.4]
  assign entriesToCheck_2_2 = _T_12870 & checkBits_2; // @[LoadQueue.scala 141:26:@11627.4]
  assign _T_12872 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11628.4]
  assign entriesToCheck_2_3 = _T_12872 & checkBits_2; // @[LoadQueue.scala 141:26:@11629.4]
  assign _T_12874 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11630.4]
  assign entriesToCheck_2_4 = _T_12874 & checkBits_2; // @[LoadQueue.scala 141:26:@11631.4]
  assign _T_12876 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11632.4]
  assign entriesToCheck_2_5 = _T_12876 & checkBits_2; // @[LoadQueue.scala 141:26:@11633.4]
  assign _T_12878 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11634.4]
  assign entriesToCheck_2_6 = _T_12878 & checkBits_2; // @[LoadQueue.scala 141:26:@11635.4]
  assign _T_12880 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11636.4]
  assign entriesToCheck_2_7 = _T_12880 & checkBits_2; // @[LoadQueue.scala 141:26:@11637.4]
  assign _T_12882 = storesToCheck_2_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11638.4]
  assign entriesToCheck_2_8 = _T_12882 & checkBits_2; // @[LoadQueue.scala 141:26:@11639.4]
  assign _T_12884 = storesToCheck_2_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11640.4]
  assign entriesToCheck_2_9 = _T_12884 & checkBits_2; // @[LoadQueue.scala 141:26:@11641.4]
  assign _T_12886 = storesToCheck_2_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11642.4]
  assign entriesToCheck_2_10 = _T_12886 & checkBits_2; // @[LoadQueue.scala 141:26:@11643.4]
  assign _T_12888 = storesToCheck_2_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11644.4]
  assign entriesToCheck_2_11 = _T_12888 & checkBits_2; // @[LoadQueue.scala 141:26:@11645.4]
  assign _T_12890 = storesToCheck_2_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11646.4]
  assign entriesToCheck_2_12 = _T_12890 & checkBits_2; // @[LoadQueue.scala 141:26:@11647.4]
  assign _T_12892 = storesToCheck_2_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11648.4]
  assign entriesToCheck_2_13 = _T_12892 & checkBits_2; // @[LoadQueue.scala 141:26:@11649.4]
  assign _T_12894 = storesToCheck_2_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11650.4]
  assign entriesToCheck_2_14 = _T_12894 & checkBits_2; // @[LoadQueue.scala 141:26:@11651.4]
  assign _T_12896 = storesToCheck_2_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11652.4]
  assign entriesToCheck_2_15 = _T_12896 & checkBits_2; // @[LoadQueue.scala 141:26:@11653.4]
  assign _T_12898 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11670.4]
  assign entriesToCheck_3_0 = _T_12898 & checkBits_3; // @[LoadQueue.scala 141:26:@11671.4]
  assign _T_12900 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11672.4]
  assign entriesToCheck_3_1 = _T_12900 & checkBits_3; // @[LoadQueue.scala 141:26:@11673.4]
  assign _T_12902 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11674.4]
  assign entriesToCheck_3_2 = _T_12902 & checkBits_3; // @[LoadQueue.scala 141:26:@11675.4]
  assign _T_12904 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11676.4]
  assign entriesToCheck_3_3 = _T_12904 & checkBits_3; // @[LoadQueue.scala 141:26:@11677.4]
  assign _T_12906 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11678.4]
  assign entriesToCheck_3_4 = _T_12906 & checkBits_3; // @[LoadQueue.scala 141:26:@11679.4]
  assign _T_12908 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11680.4]
  assign entriesToCheck_3_5 = _T_12908 & checkBits_3; // @[LoadQueue.scala 141:26:@11681.4]
  assign _T_12910 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11682.4]
  assign entriesToCheck_3_6 = _T_12910 & checkBits_3; // @[LoadQueue.scala 141:26:@11683.4]
  assign _T_12912 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11684.4]
  assign entriesToCheck_3_7 = _T_12912 & checkBits_3; // @[LoadQueue.scala 141:26:@11685.4]
  assign _T_12914 = storesToCheck_3_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11686.4]
  assign entriesToCheck_3_8 = _T_12914 & checkBits_3; // @[LoadQueue.scala 141:26:@11687.4]
  assign _T_12916 = storesToCheck_3_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11688.4]
  assign entriesToCheck_3_9 = _T_12916 & checkBits_3; // @[LoadQueue.scala 141:26:@11689.4]
  assign _T_12918 = storesToCheck_3_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11690.4]
  assign entriesToCheck_3_10 = _T_12918 & checkBits_3; // @[LoadQueue.scala 141:26:@11691.4]
  assign _T_12920 = storesToCheck_3_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11692.4]
  assign entriesToCheck_3_11 = _T_12920 & checkBits_3; // @[LoadQueue.scala 141:26:@11693.4]
  assign _T_12922 = storesToCheck_3_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11694.4]
  assign entriesToCheck_3_12 = _T_12922 & checkBits_3; // @[LoadQueue.scala 141:26:@11695.4]
  assign _T_12924 = storesToCheck_3_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11696.4]
  assign entriesToCheck_3_13 = _T_12924 & checkBits_3; // @[LoadQueue.scala 141:26:@11697.4]
  assign _T_12926 = storesToCheck_3_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11698.4]
  assign entriesToCheck_3_14 = _T_12926 & checkBits_3; // @[LoadQueue.scala 141:26:@11699.4]
  assign _T_12928 = storesToCheck_3_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11700.4]
  assign entriesToCheck_3_15 = _T_12928 & checkBits_3; // @[LoadQueue.scala 141:26:@11701.4]
  assign _T_12930 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11718.4]
  assign entriesToCheck_4_0 = _T_12930 & checkBits_4; // @[LoadQueue.scala 141:26:@11719.4]
  assign _T_12932 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11720.4]
  assign entriesToCheck_4_1 = _T_12932 & checkBits_4; // @[LoadQueue.scala 141:26:@11721.4]
  assign _T_12934 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11722.4]
  assign entriesToCheck_4_2 = _T_12934 & checkBits_4; // @[LoadQueue.scala 141:26:@11723.4]
  assign _T_12936 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11724.4]
  assign entriesToCheck_4_3 = _T_12936 & checkBits_4; // @[LoadQueue.scala 141:26:@11725.4]
  assign _T_12938 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11726.4]
  assign entriesToCheck_4_4 = _T_12938 & checkBits_4; // @[LoadQueue.scala 141:26:@11727.4]
  assign _T_12940 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11728.4]
  assign entriesToCheck_4_5 = _T_12940 & checkBits_4; // @[LoadQueue.scala 141:26:@11729.4]
  assign _T_12942 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11730.4]
  assign entriesToCheck_4_6 = _T_12942 & checkBits_4; // @[LoadQueue.scala 141:26:@11731.4]
  assign _T_12944 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11732.4]
  assign entriesToCheck_4_7 = _T_12944 & checkBits_4; // @[LoadQueue.scala 141:26:@11733.4]
  assign _T_12946 = storesToCheck_4_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11734.4]
  assign entriesToCheck_4_8 = _T_12946 & checkBits_4; // @[LoadQueue.scala 141:26:@11735.4]
  assign _T_12948 = storesToCheck_4_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11736.4]
  assign entriesToCheck_4_9 = _T_12948 & checkBits_4; // @[LoadQueue.scala 141:26:@11737.4]
  assign _T_12950 = storesToCheck_4_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11738.4]
  assign entriesToCheck_4_10 = _T_12950 & checkBits_4; // @[LoadQueue.scala 141:26:@11739.4]
  assign _T_12952 = storesToCheck_4_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11740.4]
  assign entriesToCheck_4_11 = _T_12952 & checkBits_4; // @[LoadQueue.scala 141:26:@11741.4]
  assign _T_12954 = storesToCheck_4_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11742.4]
  assign entriesToCheck_4_12 = _T_12954 & checkBits_4; // @[LoadQueue.scala 141:26:@11743.4]
  assign _T_12956 = storesToCheck_4_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11744.4]
  assign entriesToCheck_4_13 = _T_12956 & checkBits_4; // @[LoadQueue.scala 141:26:@11745.4]
  assign _T_12958 = storesToCheck_4_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11746.4]
  assign entriesToCheck_4_14 = _T_12958 & checkBits_4; // @[LoadQueue.scala 141:26:@11747.4]
  assign _T_12960 = storesToCheck_4_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11748.4]
  assign entriesToCheck_4_15 = _T_12960 & checkBits_4; // @[LoadQueue.scala 141:26:@11749.4]
  assign _T_12962 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11766.4]
  assign entriesToCheck_5_0 = _T_12962 & checkBits_5; // @[LoadQueue.scala 141:26:@11767.4]
  assign _T_12964 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11768.4]
  assign entriesToCheck_5_1 = _T_12964 & checkBits_5; // @[LoadQueue.scala 141:26:@11769.4]
  assign _T_12966 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11770.4]
  assign entriesToCheck_5_2 = _T_12966 & checkBits_5; // @[LoadQueue.scala 141:26:@11771.4]
  assign _T_12968 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11772.4]
  assign entriesToCheck_5_3 = _T_12968 & checkBits_5; // @[LoadQueue.scala 141:26:@11773.4]
  assign _T_12970 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11774.4]
  assign entriesToCheck_5_4 = _T_12970 & checkBits_5; // @[LoadQueue.scala 141:26:@11775.4]
  assign _T_12972 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11776.4]
  assign entriesToCheck_5_5 = _T_12972 & checkBits_5; // @[LoadQueue.scala 141:26:@11777.4]
  assign _T_12974 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11778.4]
  assign entriesToCheck_5_6 = _T_12974 & checkBits_5; // @[LoadQueue.scala 141:26:@11779.4]
  assign _T_12976 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11780.4]
  assign entriesToCheck_5_7 = _T_12976 & checkBits_5; // @[LoadQueue.scala 141:26:@11781.4]
  assign _T_12978 = storesToCheck_5_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11782.4]
  assign entriesToCheck_5_8 = _T_12978 & checkBits_5; // @[LoadQueue.scala 141:26:@11783.4]
  assign _T_12980 = storesToCheck_5_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11784.4]
  assign entriesToCheck_5_9 = _T_12980 & checkBits_5; // @[LoadQueue.scala 141:26:@11785.4]
  assign _T_12982 = storesToCheck_5_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11786.4]
  assign entriesToCheck_5_10 = _T_12982 & checkBits_5; // @[LoadQueue.scala 141:26:@11787.4]
  assign _T_12984 = storesToCheck_5_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11788.4]
  assign entriesToCheck_5_11 = _T_12984 & checkBits_5; // @[LoadQueue.scala 141:26:@11789.4]
  assign _T_12986 = storesToCheck_5_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11790.4]
  assign entriesToCheck_5_12 = _T_12986 & checkBits_5; // @[LoadQueue.scala 141:26:@11791.4]
  assign _T_12988 = storesToCheck_5_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11792.4]
  assign entriesToCheck_5_13 = _T_12988 & checkBits_5; // @[LoadQueue.scala 141:26:@11793.4]
  assign _T_12990 = storesToCheck_5_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11794.4]
  assign entriesToCheck_5_14 = _T_12990 & checkBits_5; // @[LoadQueue.scala 141:26:@11795.4]
  assign _T_12992 = storesToCheck_5_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11796.4]
  assign entriesToCheck_5_15 = _T_12992 & checkBits_5; // @[LoadQueue.scala 141:26:@11797.4]
  assign _T_12994 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11814.4]
  assign entriesToCheck_6_0 = _T_12994 & checkBits_6; // @[LoadQueue.scala 141:26:@11815.4]
  assign _T_12996 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11816.4]
  assign entriesToCheck_6_1 = _T_12996 & checkBits_6; // @[LoadQueue.scala 141:26:@11817.4]
  assign _T_12998 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11818.4]
  assign entriesToCheck_6_2 = _T_12998 & checkBits_6; // @[LoadQueue.scala 141:26:@11819.4]
  assign _T_13000 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11820.4]
  assign entriesToCheck_6_3 = _T_13000 & checkBits_6; // @[LoadQueue.scala 141:26:@11821.4]
  assign _T_13002 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11822.4]
  assign entriesToCheck_6_4 = _T_13002 & checkBits_6; // @[LoadQueue.scala 141:26:@11823.4]
  assign _T_13004 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11824.4]
  assign entriesToCheck_6_5 = _T_13004 & checkBits_6; // @[LoadQueue.scala 141:26:@11825.4]
  assign _T_13006 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11826.4]
  assign entriesToCheck_6_6 = _T_13006 & checkBits_6; // @[LoadQueue.scala 141:26:@11827.4]
  assign _T_13008 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11828.4]
  assign entriesToCheck_6_7 = _T_13008 & checkBits_6; // @[LoadQueue.scala 141:26:@11829.4]
  assign _T_13010 = storesToCheck_6_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11830.4]
  assign entriesToCheck_6_8 = _T_13010 & checkBits_6; // @[LoadQueue.scala 141:26:@11831.4]
  assign _T_13012 = storesToCheck_6_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11832.4]
  assign entriesToCheck_6_9 = _T_13012 & checkBits_6; // @[LoadQueue.scala 141:26:@11833.4]
  assign _T_13014 = storesToCheck_6_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11834.4]
  assign entriesToCheck_6_10 = _T_13014 & checkBits_6; // @[LoadQueue.scala 141:26:@11835.4]
  assign _T_13016 = storesToCheck_6_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11836.4]
  assign entriesToCheck_6_11 = _T_13016 & checkBits_6; // @[LoadQueue.scala 141:26:@11837.4]
  assign _T_13018 = storesToCheck_6_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11838.4]
  assign entriesToCheck_6_12 = _T_13018 & checkBits_6; // @[LoadQueue.scala 141:26:@11839.4]
  assign _T_13020 = storesToCheck_6_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11840.4]
  assign entriesToCheck_6_13 = _T_13020 & checkBits_6; // @[LoadQueue.scala 141:26:@11841.4]
  assign _T_13022 = storesToCheck_6_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11842.4]
  assign entriesToCheck_6_14 = _T_13022 & checkBits_6; // @[LoadQueue.scala 141:26:@11843.4]
  assign _T_13024 = storesToCheck_6_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11844.4]
  assign entriesToCheck_6_15 = _T_13024 & checkBits_6; // @[LoadQueue.scala 141:26:@11845.4]
  assign _T_13026 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11862.4]
  assign entriesToCheck_7_0 = _T_13026 & checkBits_7; // @[LoadQueue.scala 141:26:@11863.4]
  assign _T_13028 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11864.4]
  assign entriesToCheck_7_1 = _T_13028 & checkBits_7; // @[LoadQueue.scala 141:26:@11865.4]
  assign _T_13030 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11866.4]
  assign entriesToCheck_7_2 = _T_13030 & checkBits_7; // @[LoadQueue.scala 141:26:@11867.4]
  assign _T_13032 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11868.4]
  assign entriesToCheck_7_3 = _T_13032 & checkBits_7; // @[LoadQueue.scala 141:26:@11869.4]
  assign _T_13034 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11870.4]
  assign entriesToCheck_7_4 = _T_13034 & checkBits_7; // @[LoadQueue.scala 141:26:@11871.4]
  assign _T_13036 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11872.4]
  assign entriesToCheck_7_5 = _T_13036 & checkBits_7; // @[LoadQueue.scala 141:26:@11873.4]
  assign _T_13038 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11874.4]
  assign entriesToCheck_7_6 = _T_13038 & checkBits_7; // @[LoadQueue.scala 141:26:@11875.4]
  assign _T_13040 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11876.4]
  assign entriesToCheck_7_7 = _T_13040 & checkBits_7; // @[LoadQueue.scala 141:26:@11877.4]
  assign _T_13042 = storesToCheck_7_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11878.4]
  assign entriesToCheck_7_8 = _T_13042 & checkBits_7; // @[LoadQueue.scala 141:26:@11879.4]
  assign _T_13044 = storesToCheck_7_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11880.4]
  assign entriesToCheck_7_9 = _T_13044 & checkBits_7; // @[LoadQueue.scala 141:26:@11881.4]
  assign _T_13046 = storesToCheck_7_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11882.4]
  assign entriesToCheck_7_10 = _T_13046 & checkBits_7; // @[LoadQueue.scala 141:26:@11883.4]
  assign _T_13048 = storesToCheck_7_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11884.4]
  assign entriesToCheck_7_11 = _T_13048 & checkBits_7; // @[LoadQueue.scala 141:26:@11885.4]
  assign _T_13050 = storesToCheck_7_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11886.4]
  assign entriesToCheck_7_12 = _T_13050 & checkBits_7; // @[LoadQueue.scala 141:26:@11887.4]
  assign _T_13052 = storesToCheck_7_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11888.4]
  assign entriesToCheck_7_13 = _T_13052 & checkBits_7; // @[LoadQueue.scala 141:26:@11889.4]
  assign _T_13054 = storesToCheck_7_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11890.4]
  assign entriesToCheck_7_14 = _T_13054 & checkBits_7; // @[LoadQueue.scala 141:26:@11891.4]
  assign _T_13056 = storesToCheck_7_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11892.4]
  assign entriesToCheck_7_15 = _T_13056 & checkBits_7; // @[LoadQueue.scala 141:26:@11893.4]
  assign _T_13058 = storesToCheck_8_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11910.4]
  assign entriesToCheck_8_0 = _T_13058 & checkBits_8; // @[LoadQueue.scala 141:26:@11911.4]
  assign _T_13060 = storesToCheck_8_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11912.4]
  assign entriesToCheck_8_1 = _T_13060 & checkBits_8; // @[LoadQueue.scala 141:26:@11913.4]
  assign _T_13062 = storesToCheck_8_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11914.4]
  assign entriesToCheck_8_2 = _T_13062 & checkBits_8; // @[LoadQueue.scala 141:26:@11915.4]
  assign _T_13064 = storesToCheck_8_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11916.4]
  assign entriesToCheck_8_3 = _T_13064 & checkBits_8; // @[LoadQueue.scala 141:26:@11917.4]
  assign _T_13066 = storesToCheck_8_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11918.4]
  assign entriesToCheck_8_4 = _T_13066 & checkBits_8; // @[LoadQueue.scala 141:26:@11919.4]
  assign _T_13068 = storesToCheck_8_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11920.4]
  assign entriesToCheck_8_5 = _T_13068 & checkBits_8; // @[LoadQueue.scala 141:26:@11921.4]
  assign _T_13070 = storesToCheck_8_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11922.4]
  assign entriesToCheck_8_6 = _T_13070 & checkBits_8; // @[LoadQueue.scala 141:26:@11923.4]
  assign _T_13072 = storesToCheck_8_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11924.4]
  assign entriesToCheck_8_7 = _T_13072 & checkBits_8; // @[LoadQueue.scala 141:26:@11925.4]
  assign _T_13074 = storesToCheck_8_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11926.4]
  assign entriesToCheck_8_8 = _T_13074 & checkBits_8; // @[LoadQueue.scala 141:26:@11927.4]
  assign _T_13076 = storesToCheck_8_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11928.4]
  assign entriesToCheck_8_9 = _T_13076 & checkBits_8; // @[LoadQueue.scala 141:26:@11929.4]
  assign _T_13078 = storesToCheck_8_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11930.4]
  assign entriesToCheck_8_10 = _T_13078 & checkBits_8; // @[LoadQueue.scala 141:26:@11931.4]
  assign _T_13080 = storesToCheck_8_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11932.4]
  assign entriesToCheck_8_11 = _T_13080 & checkBits_8; // @[LoadQueue.scala 141:26:@11933.4]
  assign _T_13082 = storesToCheck_8_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11934.4]
  assign entriesToCheck_8_12 = _T_13082 & checkBits_8; // @[LoadQueue.scala 141:26:@11935.4]
  assign _T_13084 = storesToCheck_8_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11936.4]
  assign entriesToCheck_8_13 = _T_13084 & checkBits_8; // @[LoadQueue.scala 141:26:@11937.4]
  assign _T_13086 = storesToCheck_8_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11938.4]
  assign entriesToCheck_8_14 = _T_13086 & checkBits_8; // @[LoadQueue.scala 141:26:@11939.4]
  assign _T_13088 = storesToCheck_8_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11940.4]
  assign entriesToCheck_8_15 = _T_13088 & checkBits_8; // @[LoadQueue.scala 141:26:@11941.4]
  assign _T_13090 = storesToCheck_9_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@11958.4]
  assign entriesToCheck_9_0 = _T_13090 & checkBits_9; // @[LoadQueue.scala 141:26:@11959.4]
  assign _T_13092 = storesToCheck_9_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@11960.4]
  assign entriesToCheck_9_1 = _T_13092 & checkBits_9; // @[LoadQueue.scala 141:26:@11961.4]
  assign _T_13094 = storesToCheck_9_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@11962.4]
  assign entriesToCheck_9_2 = _T_13094 & checkBits_9; // @[LoadQueue.scala 141:26:@11963.4]
  assign _T_13096 = storesToCheck_9_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@11964.4]
  assign entriesToCheck_9_3 = _T_13096 & checkBits_9; // @[LoadQueue.scala 141:26:@11965.4]
  assign _T_13098 = storesToCheck_9_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@11966.4]
  assign entriesToCheck_9_4 = _T_13098 & checkBits_9; // @[LoadQueue.scala 141:26:@11967.4]
  assign _T_13100 = storesToCheck_9_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@11968.4]
  assign entriesToCheck_9_5 = _T_13100 & checkBits_9; // @[LoadQueue.scala 141:26:@11969.4]
  assign _T_13102 = storesToCheck_9_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@11970.4]
  assign entriesToCheck_9_6 = _T_13102 & checkBits_9; // @[LoadQueue.scala 141:26:@11971.4]
  assign _T_13104 = storesToCheck_9_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@11972.4]
  assign entriesToCheck_9_7 = _T_13104 & checkBits_9; // @[LoadQueue.scala 141:26:@11973.4]
  assign _T_13106 = storesToCheck_9_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@11974.4]
  assign entriesToCheck_9_8 = _T_13106 & checkBits_9; // @[LoadQueue.scala 141:26:@11975.4]
  assign _T_13108 = storesToCheck_9_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@11976.4]
  assign entriesToCheck_9_9 = _T_13108 & checkBits_9; // @[LoadQueue.scala 141:26:@11977.4]
  assign _T_13110 = storesToCheck_9_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@11978.4]
  assign entriesToCheck_9_10 = _T_13110 & checkBits_9; // @[LoadQueue.scala 141:26:@11979.4]
  assign _T_13112 = storesToCheck_9_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@11980.4]
  assign entriesToCheck_9_11 = _T_13112 & checkBits_9; // @[LoadQueue.scala 141:26:@11981.4]
  assign _T_13114 = storesToCheck_9_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@11982.4]
  assign entriesToCheck_9_12 = _T_13114 & checkBits_9; // @[LoadQueue.scala 141:26:@11983.4]
  assign _T_13116 = storesToCheck_9_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@11984.4]
  assign entriesToCheck_9_13 = _T_13116 & checkBits_9; // @[LoadQueue.scala 141:26:@11985.4]
  assign _T_13118 = storesToCheck_9_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@11986.4]
  assign entriesToCheck_9_14 = _T_13118 & checkBits_9; // @[LoadQueue.scala 141:26:@11987.4]
  assign _T_13120 = storesToCheck_9_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@11988.4]
  assign entriesToCheck_9_15 = _T_13120 & checkBits_9; // @[LoadQueue.scala 141:26:@11989.4]
  assign _T_13122 = storesToCheck_10_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12006.4]
  assign entriesToCheck_10_0 = _T_13122 & checkBits_10; // @[LoadQueue.scala 141:26:@12007.4]
  assign _T_13124 = storesToCheck_10_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12008.4]
  assign entriesToCheck_10_1 = _T_13124 & checkBits_10; // @[LoadQueue.scala 141:26:@12009.4]
  assign _T_13126 = storesToCheck_10_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12010.4]
  assign entriesToCheck_10_2 = _T_13126 & checkBits_10; // @[LoadQueue.scala 141:26:@12011.4]
  assign _T_13128 = storesToCheck_10_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12012.4]
  assign entriesToCheck_10_3 = _T_13128 & checkBits_10; // @[LoadQueue.scala 141:26:@12013.4]
  assign _T_13130 = storesToCheck_10_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12014.4]
  assign entriesToCheck_10_4 = _T_13130 & checkBits_10; // @[LoadQueue.scala 141:26:@12015.4]
  assign _T_13132 = storesToCheck_10_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12016.4]
  assign entriesToCheck_10_5 = _T_13132 & checkBits_10; // @[LoadQueue.scala 141:26:@12017.4]
  assign _T_13134 = storesToCheck_10_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12018.4]
  assign entriesToCheck_10_6 = _T_13134 & checkBits_10; // @[LoadQueue.scala 141:26:@12019.4]
  assign _T_13136 = storesToCheck_10_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12020.4]
  assign entriesToCheck_10_7 = _T_13136 & checkBits_10; // @[LoadQueue.scala 141:26:@12021.4]
  assign _T_13138 = storesToCheck_10_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12022.4]
  assign entriesToCheck_10_8 = _T_13138 & checkBits_10; // @[LoadQueue.scala 141:26:@12023.4]
  assign _T_13140 = storesToCheck_10_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12024.4]
  assign entriesToCheck_10_9 = _T_13140 & checkBits_10; // @[LoadQueue.scala 141:26:@12025.4]
  assign _T_13142 = storesToCheck_10_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12026.4]
  assign entriesToCheck_10_10 = _T_13142 & checkBits_10; // @[LoadQueue.scala 141:26:@12027.4]
  assign _T_13144 = storesToCheck_10_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12028.4]
  assign entriesToCheck_10_11 = _T_13144 & checkBits_10; // @[LoadQueue.scala 141:26:@12029.4]
  assign _T_13146 = storesToCheck_10_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12030.4]
  assign entriesToCheck_10_12 = _T_13146 & checkBits_10; // @[LoadQueue.scala 141:26:@12031.4]
  assign _T_13148 = storesToCheck_10_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12032.4]
  assign entriesToCheck_10_13 = _T_13148 & checkBits_10; // @[LoadQueue.scala 141:26:@12033.4]
  assign _T_13150 = storesToCheck_10_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12034.4]
  assign entriesToCheck_10_14 = _T_13150 & checkBits_10; // @[LoadQueue.scala 141:26:@12035.4]
  assign _T_13152 = storesToCheck_10_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12036.4]
  assign entriesToCheck_10_15 = _T_13152 & checkBits_10; // @[LoadQueue.scala 141:26:@12037.4]
  assign _T_13154 = storesToCheck_11_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12054.4]
  assign entriesToCheck_11_0 = _T_13154 & checkBits_11; // @[LoadQueue.scala 141:26:@12055.4]
  assign _T_13156 = storesToCheck_11_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12056.4]
  assign entriesToCheck_11_1 = _T_13156 & checkBits_11; // @[LoadQueue.scala 141:26:@12057.4]
  assign _T_13158 = storesToCheck_11_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12058.4]
  assign entriesToCheck_11_2 = _T_13158 & checkBits_11; // @[LoadQueue.scala 141:26:@12059.4]
  assign _T_13160 = storesToCheck_11_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12060.4]
  assign entriesToCheck_11_3 = _T_13160 & checkBits_11; // @[LoadQueue.scala 141:26:@12061.4]
  assign _T_13162 = storesToCheck_11_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12062.4]
  assign entriesToCheck_11_4 = _T_13162 & checkBits_11; // @[LoadQueue.scala 141:26:@12063.4]
  assign _T_13164 = storesToCheck_11_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12064.4]
  assign entriesToCheck_11_5 = _T_13164 & checkBits_11; // @[LoadQueue.scala 141:26:@12065.4]
  assign _T_13166 = storesToCheck_11_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12066.4]
  assign entriesToCheck_11_6 = _T_13166 & checkBits_11; // @[LoadQueue.scala 141:26:@12067.4]
  assign _T_13168 = storesToCheck_11_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12068.4]
  assign entriesToCheck_11_7 = _T_13168 & checkBits_11; // @[LoadQueue.scala 141:26:@12069.4]
  assign _T_13170 = storesToCheck_11_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12070.4]
  assign entriesToCheck_11_8 = _T_13170 & checkBits_11; // @[LoadQueue.scala 141:26:@12071.4]
  assign _T_13172 = storesToCheck_11_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12072.4]
  assign entriesToCheck_11_9 = _T_13172 & checkBits_11; // @[LoadQueue.scala 141:26:@12073.4]
  assign _T_13174 = storesToCheck_11_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12074.4]
  assign entriesToCheck_11_10 = _T_13174 & checkBits_11; // @[LoadQueue.scala 141:26:@12075.4]
  assign _T_13176 = storesToCheck_11_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12076.4]
  assign entriesToCheck_11_11 = _T_13176 & checkBits_11; // @[LoadQueue.scala 141:26:@12077.4]
  assign _T_13178 = storesToCheck_11_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12078.4]
  assign entriesToCheck_11_12 = _T_13178 & checkBits_11; // @[LoadQueue.scala 141:26:@12079.4]
  assign _T_13180 = storesToCheck_11_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12080.4]
  assign entriesToCheck_11_13 = _T_13180 & checkBits_11; // @[LoadQueue.scala 141:26:@12081.4]
  assign _T_13182 = storesToCheck_11_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12082.4]
  assign entriesToCheck_11_14 = _T_13182 & checkBits_11; // @[LoadQueue.scala 141:26:@12083.4]
  assign _T_13184 = storesToCheck_11_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12084.4]
  assign entriesToCheck_11_15 = _T_13184 & checkBits_11; // @[LoadQueue.scala 141:26:@12085.4]
  assign _T_13186 = storesToCheck_12_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12102.4]
  assign entriesToCheck_12_0 = _T_13186 & checkBits_12; // @[LoadQueue.scala 141:26:@12103.4]
  assign _T_13188 = storesToCheck_12_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12104.4]
  assign entriesToCheck_12_1 = _T_13188 & checkBits_12; // @[LoadQueue.scala 141:26:@12105.4]
  assign _T_13190 = storesToCheck_12_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12106.4]
  assign entriesToCheck_12_2 = _T_13190 & checkBits_12; // @[LoadQueue.scala 141:26:@12107.4]
  assign _T_13192 = storesToCheck_12_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12108.4]
  assign entriesToCheck_12_3 = _T_13192 & checkBits_12; // @[LoadQueue.scala 141:26:@12109.4]
  assign _T_13194 = storesToCheck_12_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12110.4]
  assign entriesToCheck_12_4 = _T_13194 & checkBits_12; // @[LoadQueue.scala 141:26:@12111.4]
  assign _T_13196 = storesToCheck_12_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12112.4]
  assign entriesToCheck_12_5 = _T_13196 & checkBits_12; // @[LoadQueue.scala 141:26:@12113.4]
  assign _T_13198 = storesToCheck_12_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12114.4]
  assign entriesToCheck_12_6 = _T_13198 & checkBits_12; // @[LoadQueue.scala 141:26:@12115.4]
  assign _T_13200 = storesToCheck_12_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12116.4]
  assign entriesToCheck_12_7 = _T_13200 & checkBits_12; // @[LoadQueue.scala 141:26:@12117.4]
  assign _T_13202 = storesToCheck_12_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12118.4]
  assign entriesToCheck_12_8 = _T_13202 & checkBits_12; // @[LoadQueue.scala 141:26:@12119.4]
  assign _T_13204 = storesToCheck_12_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12120.4]
  assign entriesToCheck_12_9 = _T_13204 & checkBits_12; // @[LoadQueue.scala 141:26:@12121.4]
  assign _T_13206 = storesToCheck_12_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12122.4]
  assign entriesToCheck_12_10 = _T_13206 & checkBits_12; // @[LoadQueue.scala 141:26:@12123.4]
  assign _T_13208 = storesToCheck_12_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12124.4]
  assign entriesToCheck_12_11 = _T_13208 & checkBits_12; // @[LoadQueue.scala 141:26:@12125.4]
  assign _T_13210 = storesToCheck_12_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12126.4]
  assign entriesToCheck_12_12 = _T_13210 & checkBits_12; // @[LoadQueue.scala 141:26:@12127.4]
  assign _T_13212 = storesToCheck_12_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12128.4]
  assign entriesToCheck_12_13 = _T_13212 & checkBits_12; // @[LoadQueue.scala 141:26:@12129.4]
  assign _T_13214 = storesToCheck_12_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12130.4]
  assign entriesToCheck_12_14 = _T_13214 & checkBits_12; // @[LoadQueue.scala 141:26:@12131.4]
  assign _T_13216 = storesToCheck_12_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12132.4]
  assign entriesToCheck_12_15 = _T_13216 & checkBits_12; // @[LoadQueue.scala 141:26:@12133.4]
  assign _T_13218 = storesToCheck_13_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12150.4]
  assign entriesToCheck_13_0 = _T_13218 & checkBits_13; // @[LoadQueue.scala 141:26:@12151.4]
  assign _T_13220 = storesToCheck_13_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12152.4]
  assign entriesToCheck_13_1 = _T_13220 & checkBits_13; // @[LoadQueue.scala 141:26:@12153.4]
  assign _T_13222 = storesToCheck_13_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12154.4]
  assign entriesToCheck_13_2 = _T_13222 & checkBits_13; // @[LoadQueue.scala 141:26:@12155.4]
  assign _T_13224 = storesToCheck_13_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12156.4]
  assign entriesToCheck_13_3 = _T_13224 & checkBits_13; // @[LoadQueue.scala 141:26:@12157.4]
  assign _T_13226 = storesToCheck_13_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12158.4]
  assign entriesToCheck_13_4 = _T_13226 & checkBits_13; // @[LoadQueue.scala 141:26:@12159.4]
  assign _T_13228 = storesToCheck_13_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12160.4]
  assign entriesToCheck_13_5 = _T_13228 & checkBits_13; // @[LoadQueue.scala 141:26:@12161.4]
  assign _T_13230 = storesToCheck_13_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12162.4]
  assign entriesToCheck_13_6 = _T_13230 & checkBits_13; // @[LoadQueue.scala 141:26:@12163.4]
  assign _T_13232 = storesToCheck_13_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12164.4]
  assign entriesToCheck_13_7 = _T_13232 & checkBits_13; // @[LoadQueue.scala 141:26:@12165.4]
  assign _T_13234 = storesToCheck_13_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12166.4]
  assign entriesToCheck_13_8 = _T_13234 & checkBits_13; // @[LoadQueue.scala 141:26:@12167.4]
  assign _T_13236 = storesToCheck_13_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12168.4]
  assign entriesToCheck_13_9 = _T_13236 & checkBits_13; // @[LoadQueue.scala 141:26:@12169.4]
  assign _T_13238 = storesToCheck_13_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12170.4]
  assign entriesToCheck_13_10 = _T_13238 & checkBits_13; // @[LoadQueue.scala 141:26:@12171.4]
  assign _T_13240 = storesToCheck_13_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12172.4]
  assign entriesToCheck_13_11 = _T_13240 & checkBits_13; // @[LoadQueue.scala 141:26:@12173.4]
  assign _T_13242 = storesToCheck_13_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12174.4]
  assign entriesToCheck_13_12 = _T_13242 & checkBits_13; // @[LoadQueue.scala 141:26:@12175.4]
  assign _T_13244 = storesToCheck_13_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12176.4]
  assign entriesToCheck_13_13 = _T_13244 & checkBits_13; // @[LoadQueue.scala 141:26:@12177.4]
  assign _T_13246 = storesToCheck_13_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12178.4]
  assign entriesToCheck_13_14 = _T_13246 & checkBits_13; // @[LoadQueue.scala 141:26:@12179.4]
  assign _T_13248 = storesToCheck_13_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12180.4]
  assign entriesToCheck_13_15 = _T_13248 & checkBits_13; // @[LoadQueue.scala 141:26:@12181.4]
  assign _T_13250 = storesToCheck_14_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12198.4]
  assign entriesToCheck_14_0 = _T_13250 & checkBits_14; // @[LoadQueue.scala 141:26:@12199.4]
  assign _T_13252 = storesToCheck_14_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12200.4]
  assign entriesToCheck_14_1 = _T_13252 & checkBits_14; // @[LoadQueue.scala 141:26:@12201.4]
  assign _T_13254 = storesToCheck_14_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12202.4]
  assign entriesToCheck_14_2 = _T_13254 & checkBits_14; // @[LoadQueue.scala 141:26:@12203.4]
  assign _T_13256 = storesToCheck_14_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12204.4]
  assign entriesToCheck_14_3 = _T_13256 & checkBits_14; // @[LoadQueue.scala 141:26:@12205.4]
  assign _T_13258 = storesToCheck_14_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12206.4]
  assign entriesToCheck_14_4 = _T_13258 & checkBits_14; // @[LoadQueue.scala 141:26:@12207.4]
  assign _T_13260 = storesToCheck_14_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12208.4]
  assign entriesToCheck_14_5 = _T_13260 & checkBits_14; // @[LoadQueue.scala 141:26:@12209.4]
  assign _T_13262 = storesToCheck_14_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12210.4]
  assign entriesToCheck_14_6 = _T_13262 & checkBits_14; // @[LoadQueue.scala 141:26:@12211.4]
  assign _T_13264 = storesToCheck_14_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12212.4]
  assign entriesToCheck_14_7 = _T_13264 & checkBits_14; // @[LoadQueue.scala 141:26:@12213.4]
  assign _T_13266 = storesToCheck_14_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12214.4]
  assign entriesToCheck_14_8 = _T_13266 & checkBits_14; // @[LoadQueue.scala 141:26:@12215.4]
  assign _T_13268 = storesToCheck_14_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12216.4]
  assign entriesToCheck_14_9 = _T_13268 & checkBits_14; // @[LoadQueue.scala 141:26:@12217.4]
  assign _T_13270 = storesToCheck_14_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12218.4]
  assign entriesToCheck_14_10 = _T_13270 & checkBits_14; // @[LoadQueue.scala 141:26:@12219.4]
  assign _T_13272 = storesToCheck_14_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12220.4]
  assign entriesToCheck_14_11 = _T_13272 & checkBits_14; // @[LoadQueue.scala 141:26:@12221.4]
  assign _T_13274 = storesToCheck_14_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12222.4]
  assign entriesToCheck_14_12 = _T_13274 & checkBits_14; // @[LoadQueue.scala 141:26:@12223.4]
  assign _T_13276 = storesToCheck_14_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12224.4]
  assign entriesToCheck_14_13 = _T_13276 & checkBits_14; // @[LoadQueue.scala 141:26:@12225.4]
  assign _T_13278 = storesToCheck_14_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12226.4]
  assign entriesToCheck_14_14 = _T_13278 & checkBits_14; // @[LoadQueue.scala 141:26:@12227.4]
  assign _T_13280 = storesToCheck_14_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12228.4]
  assign entriesToCheck_14_15 = _T_13280 & checkBits_14; // @[LoadQueue.scala 141:26:@12229.4]
  assign _T_13282 = storesToCheck_15_0 & validEntriesInStoreQ_0; // @[LoadQueue.scala 141:18:@12246.4]
  assign entriesToCheck_15_0 = _T_13282 & checkBits_15; // @[LoadQueue.scala 141:26:@12247.4]
  assign _T_13284 = storesToCheck_15_1 & validEntriesInStoreQ_1; // @[LoadQueue.scala 141:18:@12248.4]
  assign entriesToCheck_15_1 = _T_13284 & checkBits_15; // @[LoadQueue.scala 141:26:@12249.4]
  assign _T_13286 = storesToCheck_15_2 & validEntriesInStoreQ_2; // @[LoadQueue.scala 141:18:@12250.4]
  assign entriesToCheck_15_2 = _T_13286 & checkBits_15; // @[LoadQueue.scala 141:26:@12251.4]
  assign _T_13288 = storesToCheck_15_3 & validEntriesInStoreQ_3; // @[LoadQueue.scala 141:18:@12252.4]
  assign entriesToCheck_15_3 = _T_13288 & checkBits_15; // @[LoadQueue.scala 141:26:@12253.4]
  assign _T_13290 = storesToCheck_15_4 & validEntriesInStoreQ_4; // @[LoadQueue.scala 141:18:@12254.4]
  assign entriesToCheck_15_4 = _T_13290 & checkBits_15; // @[LoadQueue.scala 141:26:@12255.4]
  assign _T_13292 = storesToCheck_15_5 & validEntriesInStoreQ_5; // @[LoadQueue.scala 141:18:@12256.4]
  assign entriesToCheck_15_5 = _T_13292 & checkBits_15; // @[LoadQueue.scala 141:26:@12257.4]
  assign _T_13294 = storesToCheck_15_6 & validEntriesInStoreQ_6; // @[LoadQueue.scala 141:18:@12258.4]
  assign entriesToCheck_15_6 = _T_13294 & checkBits_15; // @[LoadQueue.scala 141:26:@12259.4]
  assign _T_13296 = storesToCheck_15_7 & validEntriesInStoreQ_7; // @[LoadQueue.scala 141:18:@12260.4]
  assign entriesToCheck_15_7 = _T_13296 & checkBits_15; // @[LoadQueue.scala 141:26:@12261.4]
  assign _T_13298 = storesToCheck_15_8 & validEntriesInStoreQ_8; // @[LoadQueue.scala 141:18:@12262.4]
  assign entriesToCheck_15_8 = _T_13298 & checkBits_15; // @[LoadQueue.scala 141:26:@12263.4]
  assign _T_13300 = storesToCheck_15_9 & validEntriesInStoreQ_9; // @[LoadQueue.scala 141:18:@12264.4]
  assign entriesToCheck_15_9 = _T_13300 & checkBits_15; // @[LoadQueue.scala 141:26:@12265.4]
  assign _T_13302 = storesToCheck_15_10 & validEntriesInStoreQ_10; // @[LoadQueue.scala 141:18:@12266.4]
  assign entriesToCheck_15_10 = _T_13302 & checkBits_15; // @[LoadQueue.scala 141:26:@12267.4]
  assign _T_13304 = storesToCheck_15_11 & validEntriesInStoreQ_11; // @[LoadQueue.scala 141:18:@12268.4]
  assign entriesToCheck_15_11 = _T_13304 & checkBits_15; // @[LoadQueue.scala 141:26:@12269.4]
  assign _T_13306 = storesToCheck_15_12 & validEntriesInStoreQ_12; // @[LoadQueue.scala 141:18:@12270.4]
  assign entriesToCheck_15_12 = _T_13306 & checkBits_15; // @[LoadQueue.scala 141:26:@12271.4]
  assign _T_13308 = storesToCheck_15_13 & validEntriesInStoreQ_13; // @[LoadQueue.scala 141:18:@12272.4]
  assign entriesToCheck_15_13 = _T_13308 & checkBits_15; // @[LoadQueue.scala 141:26:@12273.4]
  assign _T_13310 = storesToCheck_15_14 & validEntriesInStoreQ_14; // @[LoadQueue.scala 141:18:@12274.4]
  assign entriesToCheck_15_14 = _T_13310 & checkBits_15; // @[LoadQueue.scala 141:26:@12275.4]
  assign _T_13312 = storesToCheck_15_15 & validEntriesInStoreQ_15; // @[LoadQueue.scala 141:18:@12276.4]
  assign entriesToCheck_15_15 = _T_13312 & checkBits_15; // @[LoadQueue.scala 141:26:@12277.4]
  assign _T_14544 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12295.4]
  assign _T_14545 = _T_14544 & addrKnown_0; // @[LoadQueue.scala 152:41:@12296.4]
  assign _T_14546 = addrQ_0 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12297.4]
  assign conflict_0_0 = _T_14545 & _T_14546; // @[LoadQueue.scala 152:68:@12298.4]
  assign _T_14548 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12300.4]
  assign _T_14549 = _T_14548 & addrKnown_0; // @[LoadQueue.scala 152:41:@12301.4]
  assign _T_14550 = addrQ_0 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12302.4]
  assign conflict_0_1 = _T_14549 & _T_14550; // @[LoadQueue.scala 152:68:@12303.4]
  assign _T_14552 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12305.4]
  assign _T_14553 = _T_14552 & addrKnown_0; // @[LoadQueue.scala 152:41:@12306.4]
  assign _T_14554 = addrQ_0 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12307.4]
  assign conflict_0_2 = _T_14553 & _T_14554; // @[LoadQueue.scala 152:68:@12308.4]
  assign _T_14556 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12310.4]
  assign _T_14557 = _T_14556 & addrKnown_0; // @[LoadQueue.scala 152:41:@12311.4]
  assign _T_14558 = addrQ_0 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12312.4]
  assign conflict_0_3 = _T_14557 & _T_14558; // @[LoadQueue.scala 152:68:@12313.4]
  assign _T_14560 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12315.4]
  assign _T_14561 = _T_14560 & addrKnown_0; // @[LoadQueue.scala 152:41:@12316.4]
  assign _T_14562 = addrQ_0 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12317.4]
  assign conflict_0_4 = _T_14561 & _T_14562; // @[LoadQueue.scala 152:68:@12318.4]
  assign _T_14564 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12320.4]
  assign _T_14565 = _T_14564 & addrKnown_0; // @[LoadQueue.scala 152:41:@12321.4]
  assign _T_14566 = addrQ_0 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12322.4]
  assign conflict_0_5 = _T_14565 & _T_14566; // @[LoadQueue.scala 152:68:@12323.4]
  assign _T_14568 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12325.4]
  assign _T_14569 = _T_14568 & addrKnown_0; // @[LoadQueue.scala 152:41:@12326.4]
  assign _T_14570 = addrQ_0 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12327.4]
  assign conflict_0_6 = _T_14569 & _T_14570; // @[LoadQueue.scala 152:68:@12328.4]
  assign _T_14572 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12330.4]
  assign _T_14573 = _T_14572 & addrKnown_0; // @[LoadQueue.scala 152:41:@12331.4]
  assign _T_14574 = addrQ_0 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12332.4]
  assign conflict_0_7 = _T_14573 & _T_14574; // @[LoadQueue.scala 152:68:@12333.4]
  assign _T_14576 = entriesToCheck_0_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12335.4]
  assign _T_14577 = _T_14576 & addrKnown_0; // @[LoadQueue.scala 152:41:@12336.4]
  assign _T_14578 = addrQ_0 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12337.4]
  assign conflict_0_8 = _T_14577 & _T_14578; // @[LoadQueue.scala 152:68:@12338.4]
  assign _T_14580 = entriesToCheck_0_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12340.4]
  assign _T_14581 = _T_14580 & addrKnown_0; // @[LoadQueue.scala 152:41:@12341.4]
  assign _T_14582 = addrQ_0 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12342.4]
  assign conflict_0_9 = _T_14581 & _T_14582; // @[LoadQueue.scala 152:68:@12343.4]
  assign _T_14584 = entriesToCheck_0_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12345.4]
  assign _T_14585 = _T_14584 & addrKnown_0; // @[LoadQueue.scala 152:41:@12346.4]
  assign _T_14586 = addrQ_0 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12347.4]
  assign conflict_0_10 = _T_14585 & _T_14586; // @[LoadQueue.scala 152:68:@12348.4]
  assign _T_14588 = entriesToCheck_0_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12350.4]
  assign _T_14589 = _T_14588 & addrKnown_0; // @[LoadQueue.scala 152:41:@12351.4]
  assign _T_14590 = addrQ_0 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12352.4]
  assign conflict_0_11 = _T_14589 & _T_14590; // @[LoadQueue.scala 152:68:@12353.4]
  assign _T_14592 = entriesToCheck_0_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12355.4]
  assign _T_14593 = _T_14592 & addrKnown_0; // @[LoadQueue.scala 152:41:@12356.4]
  assign _T_14594 = addrQ_0 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12357.4]
  assign conflict_0_12 = _T_14593 & _T_14594; // @[LoadQueue.scala 152:68:@12358.4]
  assign _T_14596 = entriesToCheck_0_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12360.4]
  assign _T_14597 = _T_14596 & addrKnown_0; // @[LoadQueue.scala 152:41:@12361.4]
  assign _T_14598 = addrQ_0 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12362.4]
  assign conflict_0_13 = _T_14597 & _T_14598; // @[LoadQueue.scala 152:68:@12363.4]
  assign _T_14600 = entriesToCheck_0_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12365.4]
  assign _T_14601 = _T_14600 & addrKnown_0; // @[LoadQueue.scala 152:41:@12366.4]
  assign _T_14602 = addrQ_0 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12367.4]
  assign conflict_0_14 = _T_14601 & _T_14602; // @[LoadQueue.scala 152:68:@12368.4]
  assign _T_14604 = entriesToCheck_0_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12370.4]
  assign _T_14605 = _T_14604 & addrKnown_0; // @[LoadQueue.scala 152:41:@12371.4]
  assign _T_14606 = addrQ_0 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12372.4]
  assign conflict_0_15 = _T_14605 & _T_14606; // @[LoadQueue.scala 152:68:@12373.4]
  assign _T_14608 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12375.4]
  assign _T_14609 = _T_14608 & addrKnown_1; // @[LoadQueue.scala 152:41:@12376.4]
  assign _T_14610 = addrQ_1 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12377.4]
  assign conflict_1_0 = _T_14609 & _T_14610; // @[LoadQueue.scala 152:68:@12378.4]
  assign _T_14612 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12380.4]
  assign _T_14613 = _T_14612 & addrKnown_1; // @[LoadQueue.scala 152:41:@12381.4]
  assign _T_14614 = addrQ_1 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12382.4]
  assign conflict_1_1 = _T_14613 & _T_14614; // @[LoadQueue.scala 152:68:@12383.4]
  assign _T_14616 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12385.4]
  assign _T_14617 = _T_14616 & addrKnown_1; // @[LoadQueue.scala 152:41:@12386.4]
  assign _T_14618 = addrQ_1 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12387.4]
  assign conflict_1_2 = _T_14617 & _T_14618; // @[LoadQueue.scala 152:68:@12388.4]
  assign _T_14620 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12390.4]
  assign _T_14621 = _T_14620 & addrKnown_1; // @[LoadQueue.scala 152:41:@12391.4]
  assign _T_14622 = addrQ_1 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12392.4]
  assign conflict_1_3 = _T_14621 & _T_14622; // @[LoadQueue.scala 152:68:@12393.4]
  assign _T_14624 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12395.4]
  assign _T_14625 = _T_14624 & addrKnown_1; // @[LoadQueue.scala 152:41:@12396.4]
  assign _T_14626 = addrQ_1 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12397.4]
  assign conflict_1_4 = _T_14625 & _T_14626; // @[LoadQueue.scala 152:68:@12398.4]
  assign _T_14628 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12400.4]
  assign _T_14629 = _T_14628 & addrKnown_1; // @[LoadQueue.scala 152:41:@12401.4]
  assign _T_14630 = addrQ_1 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12402.4]
  assign conflict_1_5 = _T_14629 & _T_14630; // @[LoadQueue.scala 152:68:@12403.4]
  assign _T_14632 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12405.4]
  assign _T_14633 = _T_14632 & addrKnown_1; // @[LoadQueue.scala 152:41:@12406.4]
  assign _T_14634 = addrQ_1 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12407.4]
  assign conflict_1_6 = _T_14633 & _T_14634; // @[LoadQueue.scala 152:68:@12408.4]
  assign _T_14636 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12410.4]
  assign _T_14637 = _T_14636 & addrKnown_1; // @[LoadQueue.scala 152:41:@12411.4]
  assign _T_14638 = addrQ_1 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12412.4]
  assign conflict_1_7 = _T_14637 & _T_14638; // @[LoadQueue.scala 152:68:@12413.4]
  assign _T_14640 = entriesToCheck_1_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12415.4]
  assign _T_14641 = _T_14640 & addrKnown_1; // @[LoadQueue.scala 152:41:@12416.4]
  assign _T_14642 = addrQ_1 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12417.4]
  assign conflict_1_8 = _T_14641 & _T_14642; // @[LoadQueue.scala 152:68:@12418.4]
  assign _T_14644 = entriesToCheck_1_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12420.4]
  assign _T_14645 = _T_14644 & addrKnown_1; // @[LoadQueue.scala 152:41:@12421.4]
  assign _T_14646 = addrQ_1 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12422.4]
  assign conflict_1_9 = _T_14645 & _T_14646; // @[LoadQueue.scala 152:68:@12423.4]
  assign _T_14648 = entriesToCheck_1_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12425.4]
  assign _T_14649 = _T_14648 & addrKnown_1; // @[LoadQueue.scala 152:41:@12426.4]
  assign _T_14650 = addrQ_1 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12427.4]
  assign conflict_1_10 = _T_14649 & _T_14650; // @[LoadQueue.scala 152:68:@12428.4]
  assign _T_14652 = entriesToCheck_1_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12430.4]
  assign _T_14653 = _T_14652 & addrKnown_1; // @[LoadQueue.scala 152:41:@12431.4]
  assign _T_14654 = addrQ_1 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12432.4]
  assign conflict_1_11 = _T_14653 & _T_14654; // @[LoadQueue.scala 152:68:@12433.4]
  assign _T_14656 = entriesToCheck_1_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12435.4]
  assign _T_14657 = _T_14656 & addrKnown_1; // @[LoadQueue.scala 152:41:@12436.4]
  assign _T_14658 = addrQ_1 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12437.4]
  assign conflict_1_12 = _T_14657 & _T_14658; // @[LoadQueue.scala 152:68:@12438.4]
  assign _T_14660 = entriesToCheck_1_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12440.4]
  assign _T_14661 = _T_14660 & addrKnown_1; // @[LoadQueue.scala 152:41:@12441.4]
  assign _T_14662 = addrQ_1 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12442.4]
  assign conflict_1_13 = _T_14661 & _T_14662; // @[LoadQueue.scala 152:68:@12443.4]
  assign _T_14664 = entriesToCheck_1_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12445.4]
  assign _T_14665 = _T_14664 & addrKnown_1; // @[LoadQueue.scala 152:41:@12446.4]
  assign _T_14666 = addrQ_1 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12447.4]
  assign conflict_1_14 = _T_14665 & _T_14666; // @[LoadQueue.scala 152:68:@12448.4]
  assign _T_14668 = entriesToCheck_1_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12450.4]
  assign _T_14669 = _T_14668 & addrKnown_1; // @[LoadQueue.scala 152:41:@12451.4]
  assign _T_14670 = addrQ_1 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12452.4]
  assign conflict_1_15 = _T_14669 & _T_14670; // @[LoadQueue.scala 152:68:@12453.4]
  assign _T_14672 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12455.4]
  assign _T_14673 = _T_14672 & addrKnown_2; // @[LoadQueue.scala 152:41:@12456.4]
  assign _T_14674 = addrQ_2 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12457.4]
  assign conflict_2_0 = _T_14673 & _T_14674; // @[LoadQueue.scala 152:68:@12458.4]
  assign _T_14676 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12460.4]
  assign _T_14677 = _T_14676 & addrKnown_2; // @[LoadQueue.scala 152:41:@12461.4]
  assign _T_14678 = addrQ_2 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12462.4]
  assign conflict_2_1 = _T_14677 & _T_14678; // @[LoadQueue.scala 152:68:@12463.4]
  assign _T_14680 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12465.4]
  assign _T_14681 = _T_14680 & addrKnown_2; // @[LoadQueue.scala 152:41:@12466.4]
  assign _T_14682 = addrQ_2 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12467.4]
  assign conflict_2_2 = _T_14681 & _T_14682; // @[LoadQueue.scala 152:68:@12468.4]
  assign _T_14684 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12470.4]
  assign _T_14685 = _T_14684 & addrKnown_2; // @[LoadQueue.scala 152:41:@12471.4]
  assign _T_14686 = addrQ_2 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12472.4]
  assign conflict_2_3 = _T_14685 & _T_14686; // @[LoadQueue.scala 152:68:@12473.4]
  assign _T_14688 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12475.4]
  assign _T_14689 = _T_14688 & addrKnown_2; // @[LoadQueue.scala 152:41:@12476.4]
  assign _T_14690 = addrQ_2 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12477.4]
  assign conflict_2_4 = _T_14689 & _T_14690; // @[LoadQueue.scala 152:68:@12478.4]
  assign _T_14692 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12480.4]
  assign _T_14693 = _T_14692 & addrKnown_2; // @[LoadQueue.scala 152:41:@12481.4]
  assign _T_14694 = addrQ_2 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12482.4]
  assign conflict_2_5 = _T_14693 & _T_14694; // @[LoadQueue.scala 152:68:@12483.4]
  assign _T_14696 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12485.4]
  assign _T_14697 = _T_14696 & addrKnown_2; // @[LoadQueue.scala 152:41:@12486.4]
  assign _T_14698 = addrQ_2 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12487.4]
  assign conflict_2_6 = _T_14697 & _T_14698; // @[LoadQueue.scala 152:68:@12488.4]
  assign _T_14700 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12490.4]
  assign _T_14701 = _T_14700 & addrKnown_2; // @[LoadQueue.scala 152:41:@12491.4]
  assign _T_14702 = addrQ_2 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12492.4]
  assign conflict_2_7 = _T_14701 & _T_14702; // @[LoadQueue.scala 152:68:@12493.4]
  assign _T_14704 = entriesToCheck_2_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12495.4]
  assign _T_14705 = _T_14704 & addrKnown_2; // @[LoadQueue.scala 152:41:@12496.4]
  assign _T_14706 = addrQ_2 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12497.4]
  assign conflict_2_8 = _T_14705 & _T_14706; // @[LoadQueue.scala 152:68:@12498.4]
  assign _T_14708 = entriesToCheck_2_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12500.4]
  assign _T_14709 = _T_14708 & addrKnown_2; // @[LoadQueue.scala 152:41:@12501.4]
  assign _T_14710 = addrQ_2 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12502.4]
  assign conflict_2_9 = _T_14709 & _T_14710; // @[LoadQueue.scala 152:68:@12503.4]
  assign _T_14712 = entriesToCheck_2_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12505.4]
  assign _T_14713 = _T_14712 & addrKnown_2; // @[LoadQueue.scala 152:41:@12506.4]
  assign _T_14714 = addrQ_2 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12507.4]
  assign conflict_2_10 = _T_14713 & _T_14714; // @[LoadQueue.scala 152:68:@12508.4]
  assign _T_14716 = entriesToCheck_2_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12510.4]
  assign _T_14717 = _T_14716 & addrKnown_2; // @[LoadQueue.scala 152:41:@12511.4]
  assign _T_14718 = addrQ_2 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12512.4]
  assign conflict_2_11 = _T_14717 & _T_14718; // @[LoadQueue.scala 152:68:@12513.4]
  assign _T_14720 = entriesToCheck_2_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12515.4]
  assign _T_14721 = _T_14720 & addrKnown_2; // @[LoadQueue.scala 152:41:@12516.4]
  assign _T_14722 = addrQ_2 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12517.4]
  assign conflict_2_12 = _T_14721 & _T_14722; // @[LoadQueue.scala 152:68:@12518.4]
  assign _T_14724 = entriesToCheck_2_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12520.4]
  assign _T_14725 = _T_14724 & addrKnown_2; // @[LoadQueue.scala 152:41:@12521.4]
  assign _T_14726 = addrQ_2 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12522.4]
  assign conflict_2_13 = _T_14725 & _T_14726; // @[LoadQueue.scala 152:68:@12523.4]
  assign _T_14728 = entriesToCheck_2_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12525.4]
  assign _T_14729 = _T_14728 & addrKnown_2; // @[LoadQueue.scala 152:41:@12526.4]
  assign _T_14730 = addrQ_2 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12527.4]
  assign conflict_2_14 = _T_14729 & _T_14730; // @[LoadQueue.scala 152:68:@12528.4]
  assign _T_14732 = entriesToCheck_2_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12530.4]
  assign _T_14733 = _T_14732 & addrKnown_2; // @[LoadQueue.scala 152:41:@12531.4]
  assign _T_14734 = addrQ_2 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12532.4]
  assign conflict_2_15 = _T_14733 & _T_14734; // @[LoadQueue.scala 152:68:@12533.4]
  assign _T_14736 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12535.4]
  assign _T_14737 = _T_14736 & addrKnown_3; // @[LoadQueue.scala 152:41:@12536.4]
  assign _T_14738 = addrQ_3 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12537.4]
  assign conflict_3_0 = _T_14737 & _T_14738; // @[LoadQueue.scala 152:68:@12538.4]
  assign _T_14740 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12540.4]
  assign _T_14741 = _T_14740 & addrKnown_3; // @[LoadQueue.scala 152:41:@12541.4]
  assign _T_14742 = addrQ_3 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12542.4]
  assign conflict_3_1 = _T_14741 & _T_14742; // @[LoadQueue.scala 152:68:@12543.4]
  assign _T_14744 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12545.4]
  assign _T_14745 = _T_14744 & addrKnown_3; // @[LoadQueue.scala 152:41:@12546.4]
  assign _T_14746 = addrQ_3 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12547.4]
  assign conflict_3_2 = _T_14745 & _T_14746; // @[LoadQueue.scala 152:68:@12548.4]
  assign _T_14748 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12550.4]
  assign _T_14749 = _T_14748 & addrKnown_3; // @[LoadQueue.scala 152:41:@12551.4]
  assign _T_14750 = addrQ_3 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12552.4]
  assign conflict_3_3 = _T_14749 & _T_14750; // @[LoadQueue.scala 152:68:@12553.4]
  assign _T_14752 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12555.4]
  assign _T_14753 = _T_14752 & addrKnown_3; // @[LoadQueue.scala 152:41:@12556.4]
  assign _T_14754 = addrQ_3 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12557.4]
  assign conflict_3_4 = _T_14753 & _T_14754; // @[LoadQueue.scala 152:68:@12558.4]
  assign _T_14756 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12560.4]
  assign _T_14757 = _T_14756 & addrKnown_3; // @[LoadQueue.scala 152:41:@12561.4]
  assign _T_14758 = addrQ_3 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12562.4]
  assign conflict_3_5 = _T_14757 & _T_14758; // @[LoadQueue.scala 152:68:@12563.4]
  assign _T_14760 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12565.4]
  assign _T_14761 = _T_14760 & addrKnown_3; // @[LoadQueue.scala 152:41:@12566.4]
  assign _T_14762 = addrQ_3 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12567.4]
  assign conflict_3_6 = _T_14761 & _T_14762; // @[LoadQueue.scala 152:68:@12568.4]
  assign _T_14764 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12570.4]
  assign _T_14765 = _T_14764 & addrKnown_3; // @[LoadQueue.scala 152:41:@12571.4]
  assign _T_14766 = addrQ_3 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12572.4]
  assign conflict_3_7 = _T_14765 & _T_14766; // @[LoadQueue.scala 152:68:@12573.4]
  assign _T_14768 = entriesToCheck_3_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12575.4]
  assign _T_14769 = _T_14768 & addrKnown_3; // @[LoadQueue.scala 152:41:@12576.4]
  assign _T_14770 = addrQ_3 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12577.4]
  assign conflict_3_8 = _T_14769 & _T_14770; // @[LoadQueue.scala 152:68:@12578.4]
  assign _T_14772 = entriesToCheck_3_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12580.4]
  assign _T_14773 = _T_14772 & addrKnown_3; // @[LoadQueue.scala 152:41:@12581.4]
  assign _T_14774 = addrQ_3 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12582.4]
  assign conflict_3_9 = _T_14773 & _T_14774; // @[LoadQueue.scala 152:68:@12583.4]
  assign _T_14776 = entriesToCheck_3_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12585.4]
  assign _T_14777 = _T_14776 & addrKnown_3; // @[LoadQueue.scala 152:41:@12586.4]
  assign _T_14778 = addrQ_3 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12587.4]
  assign conflict_3_10 = _T_14777 & _T_14778; // @[LoadQueue.scala 152:68:@12588.4]
  assign _T_14780 = entriesToCheck_3_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12590.4]
  assign _T_14781 = _T_14780 & addrKnown_3; // @[LoadQueue.scala 152:41:@12591.4]
  assign _T_14782 = addrQ_3 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12592.4]
  assign conflict_3_11 = _T_14781 & _T_14782; // @[LoadQueue.scala 152:68:@12593.4]
  assign _T_14784 = entriesToCheck_3_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12595.4]
  assign _T_14785 = _T_14784 & addrKnown_3; // @[LoadQueue.scala 152:41:@12596.4]
  assign _T_14786 = addrQ_3 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12597.4]
  assign conflict_3_12 = _T_14785 & _T_14786; // @[LoadQueue.scala 152:68:@12598.4]
  assign _T_14788 = entriesToCheck_3_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12600.4]
  assign _T_14789 = _T_14788 & addrKnown_3; // @[LoadQueue.scala 152:41:@12601.4]
  assign _T_14790 = addrQ_3 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12602.4]
  assign conflict_3_13 = _T_14789 & _T_14790; // @[LoadQueue.scala 152:68:@12603.4]
  assign _T_14792 = entriesToCheck_3_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12605.4]
  assign _T_14793 = _T_14792 & addrKnown_3; // @[LoadQueue.scala 152:41:@12606.4]
  assign _T_14794 = addrQ_3 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12607.4]
  assign conflict_3_14 = _T_14793 & _T_14794; // @[LoadQueue.scala 152:68:@12608.4]
  assign _T_14796 = entriesToCheck_3_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12610.4]
  assign _T_14797 = _T_14796 & addrKnown_3; // @[LoadQueue.scala 152:41:@12611.4]
  assign _T_14798 = addrQ_3 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12612.4]
  assign conflict_3_15 = _T_14797 & _T_14798; // @[LoadQueue.scala 152:68:@12613.4]
  assign _T_14800 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12615.4]
  assign _T_14801 = _T_14800 & addrKnown_4; // @[LoadQueue.scala 152:41:@12616.4]
  assign _T_14802 = addrQ_4 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12617.4]
  assign conflict_4_0 = _T_14801 & _T_14802; // @[LoadQueue.scala 152:68:@12618.4]
  assign _T_14804 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12620.4]
  assign _T_14805 = _T_14804 & addrKnown_4; // @[LoadQueue.scala 152:41:@12621.4]
  assign _T_14806 = addrQ_4 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12622.4]
  assign conflict_4_1 = _T_14805 & _T_14806; // @[LoadQueue.scala 152:68:@12623.4]
  assign _T_14808 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12625.4]
  assign _T_14809 = _T_14808 & addrKnown_4; // @[LoadQueue.scala 152:41:@12626.4]
  assign _T_14810 = addrQ_4 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12627.4]
  assign conflict_4_2 = _T_14809 & _T_14810; // @[LoadQueue.scala 152:68:@12628.4]
  assign _T_14812 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12630.4]
  assign _T_14813 = _T_14812 & addrKnown_4; // @[LoadQueue.scala 152:41:@12631.4]
  assign _T_14814 = addrQ_4 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12632.4]
  assign conflict_4_3 = _T_14813 & _T_14814; // @[LoadQueue.scala 152:68:@12633.4]
  assign _T_14816 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12635.4]
  assign _T_14817 = _T_14816 & addrKnown_4; // @[LoadQueue.scala 152:41:@12636.4]
  assign _T_14818 = addrQ_4 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12637.4]
  assign conflict_4_4 = _T_14817 & _T_14818; // @[LoadQueue.scala 152:68:@12638.4]
  assign _T_14820 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12640.4]
  assign _T_14821 = _T_14820 & addrKnown_4; // @[LoadQueue.scala 152:41:@12641.4]
  assign _T_14822 = addrQ_4 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12642.4]
  assign conflict_4_5 = _T_14821 & _T_14822; // @[LoadQueue.scala 152:68:@12643.4]
  assign _T_14824 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12645.4]
  assign _T_14825 = _T_14824 & addrKnown_4; // @[LoadQueue.scala 152:41:@12646.4]
  assign _T_14826 = addrQ_4 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12647.4]
  assign conflict_4_6 = _T_14825 & _T_14826; // @[LoadQueue.scala 152:68:@12648.4]
  assign _T_14828 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12650.4]
  assign _T_14829 = _T_14828 & addrKnown_4; // @[LoadQueue.scala 152:41:@12651.4]
  assign _T_14830 = addrQ_4 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12652.4]
  assign conflict_4_7 = _T_14829 & _T_14830; // @[LoadQueue.scala 152:68:@12653.4]
  assign _T_14832 = entriesToCheck_4_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12655.4]
  assign _T_14833 = _T_14832 & addrKnown_4; // @[LoadQueue.scala 152:41:@12656.4]
  assign _T_14834 = addrQ_4 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12657.4]
  assign conflict_4_8 = _T_14833 & _T_14834; // @[LoadQueue.scala 152:68:@12658.4]
  assign _T_14836 = entriesToCheck_4_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12660.4]
  assign _T_14837 = _T_14836 & addrKnown_4; // @[LoadQueue.scala 152:41:@12661.4]
  assign _T_14838 = addrQ_4 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12662.4]
  assign conflict_4_9 = _T_14837 & _T_14838; // @[LoadQueue.scala 152:68:@12663.4]
  assign _T_14840 = entriesToCheck_4_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12665.4]
  assign _T_14841 = _T_14840 & addrKnown_4; // @[LoadQueue.scala 152:41:@12666.4]
  assign _T_14842 = addrQ_4 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12667.4]
  assign conflict_4_10 = _T_14841 & _T_14842; // @[LoadQueue.scala 152:68:@12668.4]
  assign _T_14844 = entriesToCheck_4_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12670.4]
  assign _T_14845 = _T_14844 & addrKnown_4; // @[LoadQueue.scala 152:41:@12671.4]
  assign _T_14846 = addrQ_4 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12672.4]
  assign conflict_4_11 = _T_14845 & _T_14846; // @[LoadQueue.scala 152:68:@12673.4]
  assign _T_14848 = entriesToCheck_4_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12675.4]
  assign _T_14849 = _T_14848 & addrKnown_4; // @[LoadQueue.scala 152:41:@12676.4]
  assign _T_14850 = addrQ_4 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12677.4]
  assign conflict_4_12 = _T_14849 & _T_14850; // @[LoadQueue.scala 152:68:@12678.4]
  assign _T_14852 = entriesToCheck_4_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12680.4]
  assign _T_14853 = _T_14852 & addrKnown_4; // @[LoadQueue.scala 152:41:@12681.4]
  assign _T_14854 = addrQ_4 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12682.4]
  assign conflict_4_13 = _T_14853 & _T_14854; // @[LoadQueue.scala 152:68:@12683.4]
  assign _T_14856 = entriesToCheck_4_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12685.4]
  assign _T_14857 = _T_14856 & addrKnown_4; // @[LoadQueue.scala 152:41:@12686.4]
  assign _T_14858 = addrQ_4 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12687.4]
  assign conflict_4_14 = _T_14857 & _T_14858; // @[LoadQueue.scala 152:68:@12688.4]
  assign _T_14860 = entriesToCheck_4_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12690.4]
  assign _T_14861 = _T_14860 & addrKnown_4; // @[LoadQueue.scala 152:41:@12691.4]
  assign _T_14862 = addrQ_4 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12692.4]
  assign conflict_4_15 = _T_14861 & _T_14862; // @[LoadQueue.scala 152:68:@12693.4]
  assign _T_14864 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12695.4]
  assign _T_14865 = _T_14864 & addrKnown_5; // @[LoadQueue.scala 152:41:@12696.4]
  assign _T_14866 = addrQ_5 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12697.4]
  assign conflict_5_0 = _T_14865 & _T_14866; // @[LoadQueue.scala 152:68:@12698.4]
  assign _T_14868 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12700.4]
  assign _T_14869 = _T_14868 & addrKnown_5; // @[LoadQueue.scala 152:41:@12701.4]
  assign _T_14870 = addrQ_5 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12702.4]
  assign conflict_5_1 = _T_14869 & _T_14870; // @[LoadQueue.scala 152:68:@12703.4]
  assign _T_14872 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12705.4]
  assign _T_14873 = _T_14872 & addrKnown_5; // @[LoadQueue.scala 152:41:@12706.4]
  assign _T_14874 = addrQ_5 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12707.4]
  assign conflict_5_2 = _T_14873 & _T_14874; // @[LoadQueue.scala 152:68:@12708.4]
  assign _T_14876 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12710.4]
  assign _T_14877 = _T_14876 & addrKnown_5; // @[LoadQueue.scala 152:41:@12711.4]
  assign _T_14878 = addrQ_5 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12712.4]
  assign conflict_5_3 = _T_14877 & _T_14878; // @[LoadQueue.scala 152:68:@12713.4]
  assign _T_14880 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12715.4]
  assign _T_14881 = _T_14880 & addrKnown_5; // @[LoadQueue.scala 152:41:@12716.4]
  assign _T_14882 = addrQ_5 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12717.4]
  assign conflict_5_4 = _T_14881 & _T_14882; // @[LoadQueue.scala 152:68:@12718.4]
  assign _T_14884 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12720.4]
  assign _T_14885 = _T_14884 & addrKnown_5; // @[LoadQueue.scala 152:41:@12721.4]
  assign _T_14886 = addrQ_5 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12722.4]
  assign conflict_5_5 = _T_14885 & _T_14886; // @[LoadQueue.scala 152:68:@12723.4]
  assign _T_14888 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12725.4]
  assign _T_14889 = _T_14888 & addrKnown_5; // @[LoadQueue.scala 152:41:@12726.4]
  assign _T_14890 = addrQ_5 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12727.4]
  assign conflict_5_6 = _T_14889 & _T_14890; // @[LoadQueue.scala 152:68:@12728.4]
  assign _T_14892 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12730.4]
  assign _T_14893 = _T_14892 & addrKnown_5; // @[LoadQueue.scala 152:41:@12731.4]
  assign _T_14894 = addrQ_5 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12732.4]
  assign conflict_5_7 = _T_14893 & _T_14894; // @[LoadQueue.scala 152:68:@12733.4]
  assign _T_14896 = entriesToCheck_5_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12735.4]
  assign _T_14897 = _T_14896 & addrKnown_5; // @[LoadQueue.scala 152:41:@12736.4]
  assign _T_14898 = addrQ_5 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12737.4]
  assign conflict_5_8 = _T_14897 & _T_14898; // @[LoadQueue.scala 152:68:@12738.4]
  assign _T_14900 = entriesToCheck_5_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12740.4]
  assign _T_14901 = _T_14900 & addrKnown_5; // @[LoadQueue.scala 152:41:@12741.4]
  assign _T_14902 = addrQ_5 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12742.4]
  assign conflict_5_9 = _T_14901 & _T_14902; // @[LoadQueue.scala 152:68:@12743.4]
  assign _T_14904 = entriesToCheck_5_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12745.4]
  assign _T_14905 = _T_14904 & addrKnown_5; // @[LoadQueue.scala 152:41:@12746.4]
  assign _T_14906 = addrQ_5 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12747.4]
  assign conflict_5_10 = _T_14905 & _T_14906; // @[LoadQueue.scala 152:68:@12748.4]
  assign _T_14908 = entriesToCheck_5_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12750.4]
  assign _T_14909 = _T_14908 & addrKnown_5; // @[LoadQueue.scala 152:41:@12751.4]
  assign _T_14910 = addrQ_5 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12752.4]
  assign conflict_5_11 = _T_14909 & _T_14910; // @[LoadQueue.scala 152:68:@12753.4]
  assign _T_14912 = entriesToCheck_5_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12755.4]
  assign _T_14913 = _T_14912 & addrKnown_5; // @[LoadQueue.scala 152:41:@12756.4]
  assign _T_14914 = addrQ_5 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12757.4]
  assign conflict_5_12 = _T_14913 & _T_14914; // @[LoadQueue.scala 152:68:@12758.4]
  assign _T_14916 = entriesToCheck_5_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12760.4]
  assign _T_14917 = _T_14916 & addrKnown_5; // @[LoadQueue.scala 152:41:@12761.4]
  assign _T_14918 = addrQ_5 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12762.4]
  assign conflict_5_13 = _T_14917 & _T_14918; // @[LoadQueue.scala 152:68:@12763.4]
  assign _T_14920 = entriesToCheck_5_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12765.4]
  assign _T_14921 = _T_14920 & addrKnown_5; // @[LoadQueue.scala 152:41:@12766.4]
  assign _T_14922 = addrQ_5 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12767.4]
  assign conflict_5_14 = _T_14921 & _T_14922; // @[LoadQueue.scala 152:68:@12768.4]
  assign _T_14924 = entriesToCheck_5_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12770.4]
  assign _T_14925 = _T_14924 & addrKnown_5; // @[LoadQueue.scala 152:41:@12771.4]
  assign _T_14926 = addrQ_5 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12772.4]
  assign conflict_5_15 = _T_14925 & _T_14926; // @[LoadQueue.scala 152:68:@12773.4]
  assign _T_14928 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12775.4]
  assign _T_14929 = _T_14928 & addrKnown_6; // @[LoadQueue.scala 152:41:@12776.4]
  assign _T_14930 = addrQ_6 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12777.4]
  assign conflict_6_0 = _T_14929 & _T_14930; // @[LoadQueue.scala 152:68:@12778.4]
  assign _T_14932 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12780.4]
  assign _T_14933 = _T_14932 & addrKnown_6; // @[LoadQueue.scala 152:41:@12781.4]
  assign _T_14934 = addrQ_6 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12782.4]
  assign conflict_6_1 = _T_14933 & _T_14934; // @[LoadQueue.scala 152:68:@12783.4]
  assign _T_14936 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12785.4]
  assign _T_14937 = _T_14936 & addrKnown_6; // @[LoadQueue.scala 152:41:@12786.4]
  assign _T_14938 = addrQ_6 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12787.4]
  assign conflict_6_2 = _T_14937 & _T_14938; // @[LoadQueue.scala 152:68:@12788.4]
  assign _T_14940 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12790.4]
  assign _T_14941 = _T_14940 & addrKnown_6; // @[LoadQueue.scala 152:41:@12791.4]
  assign _T_14942 = addrQ_6 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12792.4]
  assign conflict_6_3 = _T_14941 & _T_14942; // @[LoadQueue.scala 152:68:@12793.4]
  assign _T_14944 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12795.4]
  assign _T_14945 = _T_14944 & addrKnown_6; // @[LoadQueue.scala 152:41:@12796.4]
  assign _T_14946 = addrQ_6 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12797.4]
  assign conflict_6_4 = _T_14945 & _T_14946; // @[LoadQueue.scala 152:68:@12798.4]
  assign _T_14948 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12800.4]
  assign _T_14949 = _T_14948 & addrKnown_6; // @[LoadQueue.scala 152:41:@12801.4]
  assign _T_14950 = addrQ_6 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12802.4]
  assign conflict_6_5 = _T_14949 & _T_14950; // @[LoadQueue.scala 152:68:@12803.4]
  assign _T_14952 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12805.4]
  assign _T_14953 = _T_14952 & addrKnown_6; // @[LoadQueue.scala 152:41:@12806.4]
  assign _T_14954 = addrQ_6 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12807.4]
  assign conflict_6_6 = _T_14953 & _T_14954; // @[LoadQueue.scala 152:68:@12808.4]
  assign _T_14956 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12810.4]
  assign _T_14957 = _T_14956 & addrKnown_6; // @[LoadQueue.scala 152:41:@12811.4]
  assign _T_14958 = addrQ_6 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12812.4]
  assign conflict_6_7 = _T_14957 & _T_14958; // @[LoadQueue.scala 152:68:@12813.4]
  assign _T_14960 = entriesToCheck_6_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12815.4]
  assign _T_14961 = _T_14960 & addrKnown_6; // @[LoadQueue.scala 152:41:@12816.4]
  assign _T_14962 = addrQ_6 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12817.4]
  assign conflict_6_8 = _T_14961 & _T_14962; // @[LoadQueue.scala 152:68:@12818.4]
  assign _T_14964 = entriesToCheck_6_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12820.4]
  assign _T_14965 = _T_14964 & addrKnown_6; // @[LoadQueue.scala 152:41:@12821.4]
  assign _T_14966 = addrQ_6 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12822.4]
  assign conflict_6_9 = _T_14965 & _T_14966; // @[LoadQueue.scala 152:68:@12823.4]
  assign _T_14968 = entriesToCheck_6_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12825.4]
  assign _T_14969 = _T_14968 & addrKnown_6; // @[LoadQueue.scala 152:41:@12826.4]
  assign _T_14970 = addrQ_6 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12827.4]
  assign conflict_6_10 = _T_14969 & _T_14970; // @[LoadQueue.scala 152:68:@12828.4]
  assign _T_14972 = entriesToCheck_6_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12830.4]
  assign _T_14973 = _T_14972 & addrKnown_6; // @[LoadQueue.scala 152:41:@12831.4]
  assign _T_14974 = addrQ_6 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12832.4]
  assign conflict_6_11 = _T_14973 & _T_14974; // @[LoadQueue.scala 152:68:@12833.4]
  assign _T_14976 = entriesToCheck_6_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12835.4]
  assign _T_14977 = _T_14976 & addrKnown_6; // @[LoadQueue.scala 152:41:@12836.4]
  assign _T_14978 = addrQ_6 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12837.4]
  assign conflict_6_12 = _T_14977 & _T_14978; // @[LoadQueue.scala 152:68:@12838.4]
  assign _T_14980 = entriesToCheck_6_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12840.4]
  assign _T_14981 = _T_14980 & addrKnown_6; // @[LoadQueue.scala 152:41:@12841.4]
  assign _T_14982 = addrQ_6 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12842.4]
  assign conflict_6_13 = _T_14981 & _T_14982; // @[LoadQueue.scala 152:68:@12843.4]
  assign _T_14984 = entriesToCheck_6_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12845.4]
  assign _T_14985 = _T_14984 & addrKnown_6; // @[LoadQueue.scala 152:41:@12846.4]
  assign _T_14986 = addrQ_6 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12847.4]
  assign conflict_6_14 = _T_14985 & _T_14986; // @[LoadQueue.scala 152:68:@12848.4]
  assign _T_14988 = entriesToCheck_6_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12850.4]
  assign _T_14989 = _T_14988 & addrKnown_6; // @[LoadQueue.scala 152:41:@12851.4]
  assign _T_14990 = addrQ_6 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12852.4]
  assign conflict_6_15 = _T_14989 & _T_14990; // @[LoadQueue.scala 152:68:@12853.4]
  assign _T_14992 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12855.4]
  assign _T_14993 = _T_14992 & addrKnown_7; // @[LoadQueue.scala 152:41:@12856.4]
  assign _T_14994 = addrQ_7 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12857.4]
  assign conflict_7_0 = _T_14993 & _T_14994; // @[LoadQueue.scala 152:68:@12858.4]
  assign _T_14996 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12860.4]
  assign _T_14997 = _T_14996 & addrKnown_7; // @[LoadQueue.scala 152:41:@12861.4]
  assign _T_14998 = addrQ_7 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12862.4]
  assign conflict_7_1 = _T_14997 & _T_14998; // @[LoadQueue.scala 152:68:@12863.4]
  assign _T_15000 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12865.4]
  assign _T_15001 = _T_15000 & addrKnown_7; // @[LoadQueue.scala 152:41:@12866.4]
  assign _T_15002 = addrQ_7 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12867.4]
  assign conflict_7_2 = _T_15001 & _T_15002; // @[LoadQueue.scala 152:68:@12868.4]
  assign _T_15004 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12870.4]
  assign _T_15005 = _T_15004 & addrKnown_7; // @[LoadQueue.scala 152:41:@12871.4]
  assign _T_15006 = addrQ_7 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12872.4]
  assign conflict_7_3 = _T_15005 & _T_15006; // @[LoadQueue.scala 152:68:@12873.4]
  assign _T_15008 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12875.4]
  assign _T_15009 = _T_15008 & addrKnown_7; // @[LoadQueue.scala 152:41:@12876.4]
  assign _T_15010 = addrQ_7 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12877.4]
  assign conflict_7_4 = _T_15009 & _T_15010; // @[LoadQueue.scala 152:68:@12878.4]
  assign _T_15012 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12880.4]
  assign _T_15013 = _T_15012 & addrKnown_7; // @[LoadQueue.scala 152:41:@12881.4]
  assign _T_15014 = addrQ_7 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12882.4]
  assign conflict_7_5 = _T_15013 & _T_15014; // @[LoadQueue.scala 152:68:@12883.4]
  assign _T_15016 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12885.4]
  assign _T_15017 = _T_15016 & addrKnown_7; // @[LoadQueue.scala 152:41:@12886.4]
  assign _T_15018 = addrQ_7 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12887.4]
  assign conflict_7_6 = _T_15017 & _T_15018; // @[LoadQueue.scala 152:68:@12888.4]
  assign _T_15020 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12890.4]
  assign _T_15021 = _T_15020 & addrKnown_7; // @[LoadQueue.scala 152:41:@12891.4]
  assign _T_15022 = addrQ_7 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12892.4]
  assign conflict_7_7 = _T_15021 & _T_15022; // @[LoadQueue.scala 152:68:@12893.4]
  assign _T_15024 = entriesToCheck_7_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12895.4]
  assign _T_15025 = _T_15024 & addrKnown_7; // @[LoadQueue.scala 152:41:@12896.4]
  assign _T_15026 = addrQ_7 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12897.4]
  assign conflict_7_8 = _T_15025 & _T_15026; // @[LoadQueue.scala 152:68:@12898.4]
  assign _T_15028 = entriesToCheck_7_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12900.4]
  assign _T_15029 = _T_15028 & addrKnown_7; // @[LoadQueue.scala 152:41:@12901.4]
  assign _T_15030 = addrQ_7 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12902.4]
  assign conflict_7_9 = _T_15029 & _T_15030; // @[LoadQueue.scala 152:68:@12903.4]
  assign _T_15032 = entriesToCheck_7_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12905.4]
  assign _T_15033 = _T_15032 & addrKnown_7; // @[LoadQueue.scala 152:41:@12906.4]
  assign _T_15034 = addrQ_7 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12907.4]
  assign conflict_7_10 = _T_15033 & _T_15034; // @[LoadQueue.scala 152:68:@12908.4]
  assign _T_15036 = entriesToCheck_7_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12910.4]
  assign _T_15037 = _T_15036 & addrKnown_7; // @[LoadQueue.scala 152:41:@12911.4]
  assign _T_15038 = addrQ_7 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12912.4]
  assign conflict_7_11 = _T_15037 & _T_15038; // @[LoadQueue.scala 152:68:@12913.4]
  assign _T_15040 = entriesToCheck_7_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12915.4]
  assign _T_15041 = _T_15040 & addrKnown_7; // @[LoadQueue.scala 152:41:@12916.4]
  assign _T_15042 = addrQ_7 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12917.4]
  assign conflict_7_12 = _T_15041 & _T_15042; // @[LoadQueue.scala 152:68:@12918.4]
  assign _T_15044 = entriesToCheck_7_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@12920.4]
  assign _T_15045 = _T_15044 & addrKnown_7; // @[LoadQueue.scala 152:41:@12921.4]
  assign _T_15046 = addrQ_7 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@12922.4]
  assign conflict_7_13 = _T_15045 & _T_15046; // @[LoadQueue.scala 152:68:@12923.4]
  assign _T_15048 = entriesToCheck_7_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@12925.4]
  assign _T_15049 = _T_15048 & addrKnown_7; // @[LoadQueue.scala 152:41:@12926.4]
  assign _T_15050 = addrQ_7 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@12927.4]
  assign conflict_7_14 = _T_15049 & _T_15050; // @[LoadQueue.scala 152:68:@12928.4]
  assign _T_15052 = entriesToCheck_7_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@12930.4]
  assign _T_15053 = _T_15052 & addrKnown_7; // @[LoadQueue.scala 152:41:@12931.4]
  assign _T_15054 = addrQ_7 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@12932.4]
  assign conflict_7_15 = _T_15053 & _T_15054; // @[LoadQueue.scala 152:68:@12933.4]
  assign _T_15056 = entriesToCheck_8_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@12935.4]
  assign _T_15057 = _T_15056 & addrKnown_8; // @[LoadQueue.scala 152:41:@12936.4]
  assign _T_15058 = addrQ_8 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@12937.4]
  assign conflict_8_0 = _T_15057 & _T_15058; // @[LoadQueue.scala 152:68:@12938.4]
  assign _T_15060 = entriesToCheck_8_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@12940.4]
  assign _T_15061 = _T_15060 & addrKnown_8; // @[LoadQueue.scala 152:41:@12941.4]
  assign _T_15062 = addrQ_8 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@12942.4]
  assign conflict_8_1 = _T_15061 & _T_15062; // @[LoadQueue.scala 152:68:@12943.4]
  assign _T_15064 = entriesToCheck_8_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@12945.4]
  assign _T_15065 = _T_15064 & addrKnown_8; // @[LoadQueue.scala 152:41:@12946.4]
  assign _T_15066 = addrQ_8 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@12947.4]
  assign conflict_8_2 = _T_15065 & _T_15066; // @[LoadQueue.scala 152:68:@12948.4]
  assign _T_15068 = entriesToCheck_8_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@12950.4]
  assign _T_15069 = _T_15068 & addrKnown_8; // @[LoadQueue.scala 152:41:@12951.4]
  assign _T_15070 = addrQ_8 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@12952.4]
  assign conflict_8_3 = _T_15069 & _T_15070; // @[LoadQueue.scala 152:68:@12953.4]
  assign _T_15072 = entriesToCheck_8_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@12955.4]
  assign _T_15073 = _T_15072 & addrKnown_8; // @[LoadQueue.scala 152:41:@12956.4]
  assign _T_15074 = addrQ_8 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@12957.4]
  assign conflict_8_4 = _T_15073 & _T_15074; // @[LoadQueue.scala 152:68:@12958.4]
  assign _T_15076 = entriesToCheck_8_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@12960.4]
  assign _T_15077 = _T_15076 & addrKnown_8; // @[LoadQueue.scala 152:41:@12961.4]
  assign _T_15078 = addrQ_8 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@12962.4]
  assign conflict_8_5 = _T_15077 & _T_15078; // @[LoadQueue.scala 152:68:@12963.4]
  assign _T_15080 = entriesToCheck_8_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@12965.4]
  assign _T_15081 = _T_15080 & addrKnown_8; // @[LoadQueue.scala 152:41:@12966.4]
  assign _T_15082 = addrQ_8 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@12967.4]
  assign conflict_8_6 = _T_15081 & _T_15082; // @[LoadQueue.scala 152:68:@12968.4]
  assign _T_15084 = entriesToCheck_8_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@12970.4]
  assign _T_15085 = _T_15084 & addrKnown_8; // @[LoadQueue.scala 152:41:@12971.4]
  assign _T_15086 = addrQ_8 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@12972.4]
  assign conflict_8_7 = _T_15085 & _T_15086; // @[LoadQueue.scala 152:68:@12973.4]
  assign _T_15088 = entriesToCheck_8_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@12975.4]
  assign _T_15089 = _T_15088 & addrKnown_8; // @[LoadQueue.scala 152:41:@12976.4]
  assign _T_15090 = addrQ_8 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@12977.4]
  assign conflict_8_8 = _T_15089 & _T_15090; // @[LoadQueue.scala 152:68:@12978.4]
  assign _T_15092 = entriesToCheck_8_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@12980.4]
  assign _T_15093 = _T_15092 & addrKnown_8; // @[LoadQueue.scala 152:41:@12981.4]
  assign _T_15094 = addrQ_8 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@12982.4]
  assign conflict_8_9 = _T_15093 & _T_15094; // @[LoadQueue.scala 152:68:@12983.4]
  assign _T_15096 = entriesToCheck_8_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@12985.4]
  assign _T_15097 = _T_15096 & addrKnown_8; // @[LoadQueue.scala 152:41:@12986.4]
  assign _T_15098 = addrQ_8 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@12987.4]
  assign conflict_8_10 = _T_15097 & _T_15098; // @[LoadQueue.scala 152:68:@12988.4]
  assign _T_15100 = entriesToCheck_8_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@12990.4]
  assign _T_15101 = _T_15100 & addrKnown_8; // @[LoadQueue.scala 152:41:@12991.4]
  assign _T_15102 = addrQ_8 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@12992.4]
  assign conflict_8_11 = _T_15101 & _T_15102; // @[LoadQueue.scala 152:68:@12993.4]
  assign _T_15104 = entriesToCheck_8_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@12995.4]
  assign _T_15105 = _T_15104 & addrKnown_8; // @[LoadQueue.scala 152:41:@12996.4]
  assign _T_15106 = addrQ_8 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@12997.4]
  assign conflict_8_12 = _T_15105 & _T_15106; // @[LoadQueue.scala 152:68:@12998.4]
  assign _T_15108 = entriesToCheck_8_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13000.4]
  assign _T_15109 = _T_15108 & addrKnown_8; // @[LoadQueue.scala 152:41:@13001.4]
  assign _T_15110 = addrQ_8 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13002.4]
  assign conflict_8_13 = _T_15109 & _T_15110; // @[LoadQueue.scala 152:68:@13003.4]
  assign _T_15112 = entriesToCheck_8_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13005.4]
  assign _T_15113 = _T_15112 & addrKnown_8; // @[LoadQueue.scala 152:41:@13006.4]
  assign _T_15114 = addrQ_8 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13007.4]
  assign conflict_8_14 = _T_15113 & _T_15114; // @[LoadQueue.scala 152:68:@13008.4]
  assign _T_15116 = entriesToCheck_8_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13010.4]
  assign _T_15117 = _T_15116 & addrKnown_8; // @[LoadQueue.scala 152:41:@13011.4]
  assign _T_15118 = addrQ_8 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13012.4]
  assign conflict_8_15 = _T_15117 & _T_15118; // @[LoadQueue.scala 152:68:@13013.4]
  assign _T_15120 = entriesToCheck_9_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13015.4]
  assign _T_15121 = _T_15120 & addrKnown_9; // @[LoadQueue.scala 152:41:@13016.4]
  assign _T_15122 = addrQ_9 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13017.4]
  assign conflict_9_0 = _T_15121 & _T_15122; // @[LoadQueue.scala 152:68:@13018.4]
  assign _T_15124 = entriesToCheck_9_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13020.4]
  assign _T_15125 = _T_15124 & addrKnown_9; // @[LoadQueue.scala 152:41:@13021.4]
  assign _T_15126 = addrQ_9 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13022.4]
  assign conflict_9_1 = _T_15125 & _T_15126; // @[LoadQueue.scala 152:68:@13023.4]
  assign _T_15128 = entriesToCheck_9_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13025.4]
  assign _T_15129 = _T_15128 & addrKnown_9; // @[LoadQueue.scala 152:41:@13026.4]
  assign _T_15130 = addrQ_9 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13027.4]
  assign conflict_9_2 = _T_15129 & _T_15130; // @[LoadQueue.scala 152:68:@13028.4]
  assign _T_15132 = entriesToCheck_9_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13030.4]
  assign _T_15133 = _T_15132 & addrKnown_9; // @[LoadQueue.scala 152:41:@13031.4]
  assign _T_15134 = addrQ_9 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13032.4]
  assign conflict_9_3 = _T_15133 & _T_15134; // @[LoadQueue.scala 152:68:@13033.4]
  assign _T_15136 = entriesToCheck_9_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13035.4]
  assign _T_15137 = _T_15136 & addrKnown_9; // @[LoadQueue.scala 152:41:@13036.4]
  assign _T_15138 = addrQ_9 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13037.4]
  assign conflict_9_4 = _T_15137 & _T_15138; // @[LoadQueue.scala 152:68:@13038.4]
  assign _T_15140 = entriesToCheck_9_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13040.4]
  assign _T_15141 = _T_15140 & addrKnown_9; // @[LoadQueue.scala 152:41:@13041.4]
  assign _T_15142 = addrQ_9 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13042.4]
  assign conflict_9_5 = _T_15141 & _T_15142; // @[LoadQueue.scala 152:68:@13043.4]
  assign _T_15144 = entriesToCheck_9_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13045.4]
  assign _T_15145 = _T_15144 & addrKnown_9; // @[LoadQueue.scala 152:41:@13046.4]
  assign _T_15146 = addrQ_9 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13047.4]
  assign conflict_9_6 = _T_15145 & _T_15146; // @[LoadQueue.scala 152:68:@13048.4]
  assign _T_15148 = entriesToCheck_9_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13050.4]
  assign _T_15149 = _T_15148 & addrKnown_9; // @[LoadQueue.scala 152:41:@13051.4]
  assign _T_15150 = addrQ_9 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13052.4]
  assign conflict_9_7 = _T_15149 & _T_15150; // @[LoadQueue.scala 152:68:@13053.4]
  assign _T_15152 = entriesToCheck_9_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13055.4]
  assign _T_15153 = _T_15152 & addrKnown_9; // @[LoadQueue.scala 152:41:@13056.4]
  assign _T_15154 = addrQ_9 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13057.4]
  assign conflict_9_8 = _T_15153 & _T_15154; // @[LoadQueue.scala 152:68:@13058.4]
  assign _T_15156 = entriesToCheck_9_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13060.4]
  assign _T_15157 = _T_15156 & addrKnown_9; // @[LoadQueue.scala 152:41:@13061.4]
  assign _T_15158 = addrQ_9 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13062.4]
  assign conflict_9_9 = _T_15157 & _T_15158; // @[LoadQueue.scala 152:68:@13063.4]
  assign _T_15160 = entriesToCheck_9_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13065.4]
  assign _T_15161 = _T_15160 & addrKnown_9; // @[LoadQueue.scala 152:41:@13066.4]
  assign _T_15162 = addrQ_9 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13067.4]
  assign conflict_9_10 = _T_15161 & _T_15162; // @[LoadQueue.scala 152:68:@13068.4]
  assign _T_15164 = entriesToCheck_9_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13070.4]
  assign _T_15165 = _T_15164 & addrKnown_9; // @[LoadQueue.scala 152:41:@13071.4]
  assign _T_15166 = addrQ_9 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13072.4]
  assign conflict_9_11 = _T_15165 & _T_15166; // @[LoadQueue.scala 152:68:@13073.4]
  assign _T_15168 = entriesToCheck_9_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13075.4]
  assign _T_15169 = _T_15168 & addrKnown_9; // @[LoadQueue.scala 152:41:@13076.4]
  assign _T_15170 = addrQ_9 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13077.4]
  assign conflict_9_12 = _T_15169 & _T_15170; // @[LoadQueue.scala 152:68:@13078.4]
  assign _T_15172 = entriesToCheck_9_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13080.4]
  assign _T_15173 = _T_15172 & addrKnown_9; // @[LoadQueue.scala 152:41:@13081.4]
  assign _T_15174 = addrQ_9 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13082.4]
  assign conflict_9_13 = _T_15173 & _T_15174; // @[LoadQueue.scala 152:68:@13083.4]
  assign _T_15176 = entriesToCheck_9_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13085.4]
  assign _T_15177 = _T_15176 & addrKnown_9; // @[LoadQueue.scala 152:41:@13086.4]
  assign _T_15178 = addrQ_9 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13087.4]
  assign conflict_9_14 = _T_15177 & _T_15178; // @[LoadQueue.scala 152:68:@13088.4]
  assign _T_15180 = entriesToCheck_9_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13090.4]
  assign _T_15181 = _T_15180 & addrKnown_9; // @[LoadQueue.scala 152:41:@13091.4]
  assign _T_15182 = addrQ_9 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13092.4]
  assign conflict_9_15 = _T_15181 & _T_15182; // @[LoadQueue.scala 152:68:@13093.4]
  assign _T_15184 = entriesToCheck_10_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13095.4]
  assign _T_15185 = _T_15184 & addrKnown_10; // @[LoadQueue.scala 152:41:@13096.4]
  assign _T_15186 = addrQ_10 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13097.4]
  assign conflict_10_0 = _T_15185 & _T_15186; // @[LoadQueue.scala 152:68:@13098.4]
  assign _T_15188 = entriesToCheck_10_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13100.4]
  assign _T_15189 = _T_15188 & addrKnown_10; // @[LoadQueue.scala 152:41:@13101.4]
  assign _T_15190 = addrQ_10 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13102.4]
  assign conflict_10_1 = _T_15189 & _T_15190; // @[LoadQueue.scala 152:68:@13103.4]
  assign _T_15192 = entriesToCheck_10_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13105.4]
  assign _T_15193 = _T_15192 & addrKnown_10; // @[LoadQueue.scala 152:41:@13106.4]
  assign _T_15194 = addrQ_10 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13107.4]
  assign conflict_10_2 = _T_15193 & _T_15194; // @[LoadQueue.scala 152:68:@13108.4]
  assign _T_15196 = entriesToCheck_10_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13110.4]
  assign _T_15197 = _T_15196 & addrKnown_10; // @[LoadQueue.scala 152:41:@13111.4]
  assign _T_15198 = addrQ_10 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13112.4]
  assign conflict_10_3 = _T_15197 & _T_15198; // @[LoadQueue.scala 152:68:@13113.4]
  assign _T_15200 = entriesToCheck_10_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13115.4]
  assign _T_15201 = _T_15200 & addrKnown_10; // @[LoadQueue.scala 152:41:@13116.4]
  assign _T_15202 = addrQ_10 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13117.4]
  assign conflict_10_4 = _T_15201 & _T_15202; // @[LoadQueue.scala 152:68:@13118.4]
  assign _T_15204 = entriesToCheck_10_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13120.4]
  assign _T_15205 = _T_15204 & addrKnown_10; // @[LoadQueue.scala 152:41:@13121.4]
  assign _T_15206 = addrQ_10 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13122.4]
  assign conflict_10_5 = _T_15205 & _T_15206; // @[LoadQueue.scala 152:68:@13123.4]
  assign _T_15208 = entriesToCheck_10_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13125.4]
  assign _T_15209 = _T_15208 & addrKnown_10; // @[LoadQueue.scala 152:41:@13126.4]
  assign _T_15210 = addrQ_10 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13127.4]
  assign conflict_10_6 = _T_15209 & _T_15210; // @[LoadQueue.scala 152:68:@13128.4]
  assign _T_15212 = entriesToCheck_10_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13130.4]
  assign _T_15213 = _T_15212 & addrKnown_10; // @[LoadQueue.scala 152:41:@13131.4]
  assign _T_15214 = addrQ_10 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13132.4]
  assign conflict_10_7 = _T_15213 & _T_15214; // @[LoadQueue.scala 152:68:@13133.4]
  assign _T_15216 = entriesToCheck_10_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13135.4]
  assign _T_15217 = _T_15216 & addrKnown_10; // @[LoadQueue.scala 152:41:@13136.4]
  assign _T_15218 = addrQ_10 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13137.4]
  assign conflict_10_8 = _T_15217 & _T_15218; // @[LoadQueue.scala 152:68:@13138.4]
  assign _T_15220 = entriesToCheck_10_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13140.4]
  assign _T_15221 = _T_15220 & addrKnown_10; // @[LoadQueue.scala 152:41:@13141.4]
  assign _T_15222 = addrQ_10 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13142.4]
  assign conflict_10_9 = _T_15221 & _T_15222; // @[LoadQueue.scala 152:68:@13143.4]
  assign _T_15224 = entriesToCheck_10_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13145.4]
  assign _T_15225 = _T_15224 & addrKnown_10; // @[LoadQueue.scala 152:41:@13146.4]
  assign _T_15226 = addrQ_10 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13147.4]
  assign conflict_10_10 = _T_15225 & _T_15226; // @[LoadQueue.scala 152:68:@13148.4]
  assign _T_15228 = entriesToCheck_10_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13150.4]
  assign _T_15229 = _T_15228 & addrKnown_10; // @[LoadQueue.scala 152:41:@13151.4]
  assign _T_15230 = addrQ_10 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13152.4]
  assign conflict_10_11 = _T_15229 & _T_15230; // @[LoadQueue.scala 152:68:@13153.4]
  assign _T_15232 = entriesToCheck_10_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13155.4]
  assign _T_15233 = _T_15232 & addrKnown_10; // @[LoadQueue.scala 152:41:@13156.4]
  assign _T_15234 = addrQ_10 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13157.4]
  assign conflict_10_12 = _T_15233 & _T_15234; // @[LoadQueue.scala 152:68:@13158.4]
  assign _T_15236 = entriesToCheck_10_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13160.4]
  assign _T_15237 = _T_15236 & addrKnown_10; // @[LoadQueue.scala 152:41:@13161.4]
  assign _T_15238 = addrQ_10 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13162.4]
  assign conflict_10_13 = _T_15237 & _T_15238; // @[LoadQueue.scala 152:68:@13163.4]
  assign _T_15240 = entriesToCheck_10_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13165.4]
  assign _T_15241 = _T_15240 & addrKnown_10; // @[LoadQueue.scala 152:41:@13166.4]
  assign _T_15242 = addrQ_10 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13167.4]
  assign conflict_10_14 = _T_15241 & _T_15242; // @[LoadQueue.scala 152:68:@13168.4]
  assign _T_15244 = entriesToCheck_10_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13170.4]
  assign _T_15245 = _T_15244 & addrKnown_10; // @[LoadQueue.scala 152:41:@13171.4]
  assign _T_15246 = addrQ_10 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13172.4]
  assign conflict_10_15 = _T_15245 & _T_15246; // @[LoadQueue.scala 152:68:@13173.4]
  assign _T_15248 = entriesToCheck_11_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13175.4]
  assign _T_15249 = _T_15248 & addrKnown_11; // @[LoadQueue.scala 152:41:@13176.4]
  assign _T_15250 = addrQ_11 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13177.4]
  assign conflict_11_0 = _T_15249 & _T_15250; // @[LoadQueue.scala 152:68:@13178.4]
  assign _T_15252 = entriesToCheck_11_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13180.4]
  assign _T_15253 = _T_15252 & addrKnown_11; // @[LoadQueue.scala 152:41:@13181.4]
  assign _T_15254 = addrQ_11 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13182.4]
  assign conflict_11_1 = _T_15253 & _T_15254; // @[LoadQueue.scala 152:68:@13183.4]
  assign _T_15256 = entriesToCheck_11_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13185.4]
  assign _T_15257 = _T_15256 & addrKnown_11; // @[LoadQueue.scala 152:41:@13186.4]
  assign _T_15258 = addrQ_11 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13187.4]
  assign conflict_11_2 = _T_15257 & _T_15258; // @[LoadQueue.scala 152:68:@13188.4]
  assign _T_15260 = entriesToCheck_11_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13190.4]
  assign _T_15261 = _T_15260 & addrKnown_11; // @[LoadQueue.scala 152:41:@13191.4]
  assign _T_15262 = addrQ_11 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13192.4]
  assign conflict_11_3 = _T_15261 & _T_15262; // @[LoadQueue.scala 152:68:@13193.4]
  assign _T_15264 = entriesToCheck_11_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13195.4]
  assign _T_15265 = _T_15264 & addrKnown_11; // @[LoadQueue.scala 152:41:@13196.4]
  assign _T_15266 = addrQ_11 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13197.4]
  assign conflict_11_4 = _T_15265 & _T_15266; // @[LoadQueue.scala 152:68:@13198.4]
  assign _T_15268 = entriesToCheck_11_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13200.4]
  assign _T_15269 = _T_15268 & addrKnown_11; // @[LoadQueue.scala 152:41:@13201.4]
  assign _T_15270 = addrQ_11 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13202.4]
  assign conflict_11_5 = _T_15269 & _T_15270; // @[LoadQueue.scala 152:68:@13203.4]
  assign _T_15272 = entriesToCheck_11_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13205.4]
  assign _T_15273 = _T_15272 & addrKnown_11; // @[LoadQueue.scala 152:41:@13206.4]
  assign _T_15274 = addrQ_11 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13207.4]
  assign conflict_11_6 = _T_15273 & _T_15274; // @[LoadQueue.scala 152:68:@13208.4]
  assign _T_15276 = entriesToCheck_11_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13210.4]
  assign _T_15277 = _T_15276 & addrKnown_11; // @[LoadQueue.scala 152:41:@13211.4]
  assign _T_15278 = addrQ_11 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13212.4]
  assign conflict_11_7 = _T_15277 & _T_15278; // @[LoadQueue.scala 152:68:@13213.4]
  assign _T_15280 = entriesToCheck_11_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13215.4]
  assign _T_15281 = _T_15280 & addrKnown_11; // @[LoadQueue.scala 152:41:@13216.4]
  assign _T_15282 = addrQ_11 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13217.4]
  assign conflict_11_8 = _T_15281 & _T_15282; // @[LoadQueue.scala 152:68:@13218.4]
  assign _T_15284 = entriesToCheck_11_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13220.4]
  assign _T_15285 = _T_15284 & addrKnown_11; // @[LoadQueue.scala 152:41:@13221.4]
  assign _T_15286 = addrQ_11 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13222.4]
  assign conflict_11_9 = _T_15285 & _T_15286; // @[LoadQueue.scala 152:68:@13223.4]
  assign _T_15288 = entriesToCheck_11_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13225.4]
  assign _T_15289 = _T_15288 & addrKnown_11; // @[LoadQueue.scala 152:41:@13226.4]
  assign _T_15290 = addrQ_11 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13227.4]
  assign conflict_11_10 = _T_15289 & _T_15290; // @[LoadQueue.scala 152:68:@13228.4]
  assign _T_15292 = entriesToCheck_11_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13230.4]
  assign _T_15293 = _T_15292 & addrKnown_11; // @[LoadQueue.scala 152:41:@13231.4]
  assign _T_15294 = addrQ_11 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13232.4]
  assign conflict_11_11 = _T_15293 & _T_15294; // @[LoadQueue.scala 152:68:@13233.4]
  assign _T_15296 = entriesToCheck_11_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13235.4]
  assign _T_15297 = _T_15296 & addrKnown_11; // @[LoadQueue.scala 152:41:@13236.4]
  assign _T_15298 = addrQ_11 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13237.4]
  assign conflict_11_12 = _T_15297 & _T_15298; // @[LoadQueue.scala 152:68:@13238.4]
  assign _T_15300 = entriesToCheck_11_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13240.4]
  assign _T_15301 = _T_15300 & addrKnown_11; // @[LoadQueue.scala 152:41:@13241.4]
  assign _T_15302 = addrQ_11 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13242.4]
  assign conflict_11_13 = _T_15301 & _T_15302; // @[LoadQueue.scala 152:68:@13243.4]
  assign _T_15304 = entriesToCheck_11_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13245.4]
  assign _T_15305 = _T_15304 & addrKnown_11; // @[LoadQueue.scala 152:41:@13246.4]
  assign _T_15306 = addrQ_11 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13247.4]
  assign conflict_11_14 = _T_15305 & _T_15306; // @[LoadQueue.scala 152:68:@13248.4]
  assign _T_15308 = entriesToCheck_11_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13250.4]
  assign _T_15309 = _T_15308 & addrKnown_11; // @[LoadQueue.scala 152:41:@13251.4]
  assign _T_15310 = addrQ_11 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13252.4]
  assign conflict_11_15 = _T_15309 & _T_15310; // @[LoadQueue.scala 152:68:@13253.4]
  assign _T_15312 = entriesToCheck_12_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13255.4]
  assign _T_15313 = _T_15312 & addrKnown_12; // @[LoadQueue.scala 152:41:@13256.4]
  assign _T_15314 = addrQ_12 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13257.4]
  assign conflict_12_0 = _T_15313 & _T_15314; // @[LoadQueue.scala 152:68:@13258.4]
  assign _T_15316 = entriesToCheck_12_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13260.4]
  assign _T_15317 = _T_15316 & addrKnown_12; // @[LoadQueue.scala 152:41:@13261.4]
  assign _T_15318 = addrQ_12 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13262.4]
  assign conflict_12_1 = _T_15317 & _T_15318; // @[LoadQueue.scala 152:68:@13263.4]
  assign _T_15320 = entriesToCheck_12_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13265.4]
  assign _T_15321 = _T_15320 & addrKnown_12; // @[LoadQueue.scala 152:41:@13266.4]
  assign _T_15322 = addrQ_12 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13267.4]
  assign conflict_12_2 = _T_15321 & _T_15322; // @[LoadQueue.scala 152:68:@13268.4]
  assign _T_15324 = entriesToCheck_12_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13270.4]
  assign _T_15325 = _T_15324 & addrKnown_12; // @[LoadQueue.scala 152:41:@13271.4]
  assign _T_15326 = addrQ_12 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13272.4]
  assign conflict_12_3 = _T_15325 & _T_15326; // @[LoadQueue.scala 152:68:@13273.4]
  assign _T_15328 = entriesToCheck_12_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13275.4]
  assign _T_15329 = _T_15328 & addrKnown_12; // @[LoadQueue.scala 152:41:@13276.4]
  assign _T_15330 = addrQ_12 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13277.4]
  assign conflict_12_4 = _T_15329 & _T_15330; // @[LoadQueue.scala 152:68:@13278.4]
  assign _T_15332 = entriesToCheck_12_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13280.4]
  assign _T_15333 = _T_15332 & addrKnown_12; // @[LoadQueue.scala 152:41:@13281.4]
  assign _T_15334 = addrQ_12 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13282.4]
  assign conflict_12_5 = _T_15333 & _T_15334; // @[LoadQueue.scala 152:68:@13283.4]
  assign _T_15336 = entriesToCheck_12_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13285.4]
  assign _T_15337 = _T_15336 & addrKnown_12; // @[LoadQueue.scala 152:41:@13286.4]
  assign _T_15338 = addrQ_12 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13287.4]
  assign conflict_12_6 = _T_15337 & _T_15338; // @[LoadQueue.scala 152:68:@13288.4]
  assign _T_15340 = entriesToCheck_12_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13290.4]
  assign _T_15341 = _T_15340 & addrKnown_12; // @[LoadQueue.scala 152:41:@13291.4]
  assign _T_15342 = addrQ_12 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13292.4]
  assign conflict_12_7 = _T_15341 & _T_15342; // @[LoadQueue.scala 152:68:@13293.4]
  assign _T_15344 = entriesToCheck_12_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13295.4]
  assign _T_15345 = _T_15344 & addrKnown_12; // @[LoadQueue.scala 152:41:@13296.4]
  assign _T_15346 = addrQ_12 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13297.4]
  assign conflict_12_8 = _T_15345 & _T_15346; // @[LoadQueue.scala 152:68:@13298.4]
  assign _T_15348 = entriesToCheck_12_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13300.4]
  assign _T_15349 = _T_15348 & addrKnown_12; // @[LoadQueue.scala 152:41:@13301.4]
  assign _T_15350 = addrQ_12 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13302.4]
  assign conflict_12_9 = _T_15349 & _T_15350; // @[LoadQueue.scala 152:68:@13303.4]
  assign _T_15352 = entriesToCheck_12_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13305.4]
  assign _T_15353 = _T_15352 & addrKnown_12; // @[LoadQueue.scala 152:41:@13306.4]
  assign _T_15354 = addrQ_12 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13307.4]
  assign conflict_12_10 = _T_15353 & _T_15354; // @[LoadQueue.scala 152:68:@13308.4]
  assign _T_15356 = entriesToCheck_12_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13310.4]
  assign _T_15357 = _T_15356 & addrKnown_12; // @[LoadQueue.scala 152:41:@13311.4]
  assign _T_15358 = addrQ_12 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13312.4]
  assign conflict_12_11 = _T_15357 & _T_15358; // @[LoadQueue.scala 152:68:@13313.4]
  assign _T_15360 = entriesToCheck_12_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13315.4]
  assign _T_15361 = _T_15360 & addrKnown_12; // @[LoadQueue.scala 152:41:@13316.4]
  assign _T_15362 = addrQ_12 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13317.4]
  assign conflict_12_12 = _T_15361 & _T_15362; // @[LoadQueue.scala 152:68:@13318.4]
  assign _T_15364 = entriesToCheck_12_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13320.4]
  assign _T_15365 = _T_15364 & addrKnown_12; // @[LoadQueue.scala 152:41:@13321.4]
  assign _T_15366 = addrQ_12 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13322.4]
  assign conflict_12_13 = _T_15365 & _T_15366; // @[LoadQueue.scala 152:68:@13323.4]
  assign _T_15368 = entriesToCheck_12_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13325.4]
  assign _T_15369 = _T_15368 & addrKnown_12; // @[LoadQueue.scala 152:41:@13326.4]
  assign _T_15370 = addrQ_12 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13327.4]
  assign conflict_12_14 = _T_15369 & _T_15370; // @[LoadQueue.scala 152:68:@13328.4]
  assign _T_15372 = entriesToCheck_12_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13330.4]
  assign _T_15373 = _T_15372 & addrKnown_12; // @[LoadQueue.scala 152:41:@13331.4]
  assign _T_15374 = addrQ_12 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13332.4]
  assign conflict_12_15 = _T_15373 & _T_15374; // @[LoadQueue.scala 152:68:@13333.4]
  assign _T_15376 = entriesToCheck_13_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13335.4]
  assign _T_15377 = _T_15376 & addrKnown_13; // @[LoadQueue.scala 152:41:@13336.4]
  assign _T_15378 = addrQ_13 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13337.4]
  assign conflict_13_0 = _T_15377 & _T_15378; // @[LoadQueue.scala 152:68:@13338.4]
  assign _T_15380 = entriesToCheck_13_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13340.4]
  assign _T_15381 = _T_15380 & addrKnown_13; // @[LoadQueue.scala 152:41:@13341.4]
  assign _T_15382 = addrQ_13 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13342.4]
  assign conflict_13_1 = _T_15381 & _T_15382; // @[LoadQueue.scala 152:68:@13343.4]
  assign _T_15384 = entriesToCheck_13_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13345.4]
  assign _T_15385 = _T_15384 & addrKnown_13; // @[LoadQueue.scala 152:41:@13346.4]
  assign _T_15386 = addrQ_13 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13347.4]
  assign conflict_13_2 = _T_15385 & _T_15386; // @[LoadQueue.scala 152:68:@13348.4]
  assign _T_15388 = entriesToCheck_13_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13350.4]
  assign _T_15389 = _T_15388 & addrKnown_13; // @[LoadQueue.scala 152:41:@13351.4]
  assign _T_15390 = addrQ_13 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13352.4]
  assign conflict_13_3 = _T_15389 & _T_15390; // @[LoadQueue.scala 152:68:@13353.4]
  assign _T_15392 = entriesToCheck_13_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13355.4]
  assign _T_15393 = _T_15392 & addrKnown_13; // @[LoadQueue.scala 152:41:@13356.4]
  assign _T_15394 = addrQ_13 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13357.4]
  assign conflict_13_4 = _T_15393 & _T_15394; // @[LoadQueue.scala 152:68:@13358.4]
  assign _T_15396 = entriesToCheck_13_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13360.4]
  assign _T_15397 = _T_15396 & addrKnown_13; // @[LoadQueue.scala 152:41:@13361.4]
  assign _T_15398 = addrQ_13 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13362.4]
  assign conflict_13_5 = _T_15397 & _T_15398; // @[LoadQueue.scala 152:68:@13363.4]
  assign _T_15400 = entriesToCheck_13_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13365.4]
  assign _T_15401 = _T_15400 & addrKnown_13; // @[LoadQueue.scala 152:41:@13366.4]
  assign _T_15402 = addrQ_13 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13367.4]
  assign conflict_13_6 = _T_15401 & _T_15402; // @[LoadQueue.scala 152:68:@13368.4]
  assign _T_15404 = entriesToCheck_13_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13370.4]
  assign _T_15405 = _T_15404 & addrKnown_13; // @[LoadQueue.scala 152:41:@13371.4]
  assign _T_15406 = addrQ_13 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13372.4]
  assign conflict_13_7 = _T_15405 & _T_15406; // @[LoadQueue.scala 152:68:@13373.4]
  assign _T_15408 = entriesToCheck_13_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13375.4]
  assign _T_15409 = _T_15408 & addrKnown_13; // @[LoadQueue.scala 152:41:@13376.4]
  assign _T_15410 = addrQ_13 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13377.4]
  assign conflict_13_8 = _T_15409 & _T_15410; // @[LoadQueue.scala 152:68:@13378.4]
  assign _T_15412 = entriesToCheck_13_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13380.4]
  assign _T_15413 = _T_15412 & addrKnown_13; // @[LoadQueue.scala 152:41:@13381.4]
  assign _T_15414 = addrQ_13 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13382.4]
  assign conflict_13_9 = _T_15413 & _T_15414; // @[LoadQueue.scala 152:68:@13383.4]
  assign _T_15416 = entriesToCheck_13_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13385.4]
  assign _T_15417 = _T_15416 & addrKnown_13; // @[LoadQueue.scala 152:41:@13386.4]
  assign _T_15418 = addrQ_13 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13387.4]
  assign conflict_13_10 = _T_15417 & _T_15418; // @[LoadQueue.scala 152:68:@13388.4]
  assign _T_15420 = entriesToCheck_13_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13390.4]
  assign _T_15421 = _T_15420 & addrKnown_13; // @[LoadQueue.scala 152:41:@13391.4]
  assign _T_15422 = addrQ_13 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13392.4]
  assign conflict_13_11 = _T_15421 & _T_15422; // @[LoadQueue.scala 152:68:@13393.4]
  assign _T_15424 = entriesToCheck_13_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13395.4]
  assign _T_15425 = _T_15424 & addrKnown_13; // @[LoadQueue.scala 152:41:@13396.4]
  assign _T_15426 = addrQ_13 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13397.4]
  assign conflict_13_12 = _T_15425 & _T_15426; // @[LoadQueue.scala 152:68:@13398.4]
  assign _T_15428 = entriesToCheck_13_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13400.4]
  assign _T_15429 = _T_15428 & addrKnown_13; // @[LoadQueue.scala 152:41:@13401.4]
  assign _T_15430 = addrQ_13 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13402.4]
  assign conflict_13_13 = _T_15429 & _T_15430; // @[LoadQueue.scala 152:68:@13403.4]
  assign _T_15432 = entriesToCheck_13_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13405.4]
  assign _T_15433 = _T_15432 & addrKnown_13; // @[LoadQueue.scala 152:41:@13406.4]
  assign _T_15434 = addrQ_13 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13407.4]
  assign conflict_13_14 = _T_15433 & _T_15434; // @[LoadQueue.scala 152:68:@13408.4]
  assign _T_15436 = entriesToCheck_13_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13410.4]
  assign _T_15437 = _T_15436 & addrKnown_13; // @[LoadQueue.scala 152:41:@13411.4]
  assign _T_15438 = addrQ_13 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13412.4]
  assign conflict_13_15 = _T_15437 & _T_15438; // @[LoadQueue.scala 152:68:@13413.4]
  assign _T_15440 = entriesToCheck_14_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13415.4]
  assign _T_15441 = _T_15440 & addrKnown_14; // @[LoadQueue.scala 152:41:@13416.4]
  assign _T_15442 = addrQ_14 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13417.4]
  assign conflict_14_0 = _T_15441 & _T_15442; // @[LoadQueue.scala 152:68:@13418.4]
  assign _T_15444 = entriesToCheck_14_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13420.4]
  assign _T_15445 = _T_15444 & addrKnown_14; // @[LoadQueue.scala 152:41:@13421.4]
  assign _T_15446 = addrQ_14 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13422.4]
  assign conflict_14_1 = _T_15445 & _T_15446; // @[LoadQueue.scala 152:68:@13423.4]
  assign _T_15448 = entriesToCheck_14_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13425.4]
  assign _T_15449 = _T_15448 & addrKnown_14; // @[LoadQueue.scala 152:41:@13426.4]
  assign _T_15450 = addrQ_14 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13427.4]
  assign conflict_14_2 = _T_15449 & _T_15450; // @[LoadQueue.scala 152:68:@13428.4]
  assign _T_15452 = entriesToCheck_14_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13430.4]
  assign _T_15453 = _T_15452 & addrKnown_14; // @[LoadQueue.scala 152:41:@13431.4]
  assign _T_15454 = addrQ_14 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13432.4]
  assign conflict_14_3 = _T_15453 & _T_15454; // @[LoadQueue.scala 152:68:@13433.4]
  assign _T_15456 = entriesToCheck_14_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13435.4]
  assign _T_15457 = _T_15456 & addrKnown_14; // @[LoadQueue.scala 152:41:@13436.4]
  assign _T_15458 = addrQ_14 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13437.4]
  assign conflict_14_4 = _T_15457 & _T_15458; // @[LoadQueue.scala 152:68:@13438.4]
  assign _T_15460 = entriesToCheck_14_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13440.4]
  assign _T_15461 = _T_15460 & addrKnown_14; // @[LoadQueue.scala 152:41:@13441.4]
  assign _T_15462 = addrQ_14 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13442.4]
  assign conflict_14_5 = _T_15461 & _T_15462; // @[LoadQueue.scala 152:68:@13443.4]
  assign _T_15464 = entriesToCheck_14_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13445.4]
  assign _T_15465 = _T_15464 & addrKnown_14; // @[LoadQueue.scala 152:41:@13446.4]
  assign _T_15466 = addrQ_14 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13447.4]
  assign conflict_14_6 = _T_15465 & _T_15466; // @[LoadQueue.scala 152:68:@13448.4]
  assign _T_15468 = entriesToCheck_14_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13450.4]
  assign _T_15469 = _T_15468 & addrKnown_14; // @[LoadQueue.scala 152:41:@13451.4]
  assign _T_15470 = addrQ_14 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13452.4]
  assign conflict_14_7 = _T_15469 & _T_15470; // @[LoadQueue.scala 152:68:@13453.4]
  assign _T_15472 = entriesToCheck_14_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13455.4]
  assign _T_15473 = _T_15472 & addrKnown_14; // @[LoadQueue.scala 152:41:@13456.4]
  assign _T_15474 = addrQ_14 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13457.4]
  assign conflict_14_8 = _T_15473 & _T_15474; // @[LoadQueue.scala 152:68:@13458.4]
  assign _T_15476 = entriesToCheck_14_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13460.4]
  assign _T_15477 = _T_15476 & addrKnown_14; // @[LoadQueue.scala 152:41:@13461.4]
  assign _T_15478 = addrQ_14 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13462.4]
  assign conflict_14_9 = _T_15477 & _T_15478; // @[LoadQueue.scala 152:68:@13463.4]
  assign _T_15480 = entriesToCheck_14_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13465.4]
  assign _T_15481 = _T_15480 & addrKnown_14; // @[LoadQueue.scala 152:41:@13466.4]
  assign _T_15482 = addrQ_14 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13467.4]
  assign conflict_14_10 = _T_15481 & _T_15482; // @[LoadQueue.scala 152:68:@13468.4]
  assign _T_15484 = entriesToCheck_14_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13470.4]
  assign _T_15485 = _T_15484 & addrKnown_14; // @[LoadQueue.scala 152:41:@13471.4]
  assign _T_15486 = addrQ_14 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13472.4]
  assign conflict_14_11 = _T_15485 & _T_15486; // @[LoadQueue.scala 152:68:@13473.4]
  assign _T_15488 = entriesToCheck_14_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13475.4]
  assign _T_15489 = _T_15488 & addrKnown_14; // @[LoadQueue.scala 152:41:@13476.4]
  assign _T_15490 = addrQ_14 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13477.4]
  assign conflict_14_12 = _T_15489 & _T_15490; // @[LoadQueue.scala 152:68:@13478.4]
  assign _T_15492 = entriesToCheck_14_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13480.4]
  assign _T_15493 = _T_15492 & addrKnown_14; // @[LoadQueue.scala 152:41:@13481.4]
  assign _T_15494 = addrQ_14 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13482.4]
  assign conflict_14_13 = _T_15493 & _T_15494; // @[LoadQueue.scala 152:68:@13483.4]
  assign _T_15496 = entriesToCheck_14_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13485.4]
  assign _T_15497 = _T_15496 & addrKnown_14; // @[LoadQueue.scala 152:41:@13486.4]
  assign _T_15498 = addrQ_14 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13487.4]
  assign conflict_14_14 = _T_15497 & _T_15498; // @[LoadQueue.scala 152:68:@13488.4]
  assign _T_15500 = entriesToCheck_14_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13490.4]
  assign _T_15501 = _T_15500 & addrKnown_14; // @[LoadQueue.scala 152:41:@13491.4]
  assign _T_15502 = addrQ_14 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13492.4]
  assign conflict_14_15 = _T_15501 & _T_15502; // @[LoadQueue.scala 152:68:@13493.4]
  assign _T_15504 = entriesToCheck_15_0 & io_storeAddrDone_0; // @[LoadQueue.scala 151:92:@13495.4]
  assign _T_15505 = _T_15504 & addrKnown_15; // @[LoadQueue.scala 152:41:@13496.4]
  assign _T_15506 = addrQ_15 == io_storeAddrQueue_0; // @[LoadQueue.scala 153:30:@13497.4]
  assign conflict_15_0 = _T_15505 & _T_15506; // @[LoadQueue.scala 152:68:@13498.4]
  assign _T_15508 = entriesToCheck_15_1 & io_storeAddrDone_1; // @[LoadQueue.scala 151:92:@13500.4]
  assign _T_15509 = _T_15508 & addrKnown_15; // @[LoadQueue.scala 152:41:@13501.4]
  assign _T_15510 = addrQ_15 == io_storeAddrQueue_1; // @[LoadQueue.scala 153:30:@13502.4]
  assign conflict_15_1 = _T_15509 & _T_15510; // @[LoadQueue.scala 152:68:@13503.4]
  assign _T_15512 = entriesToCheck_15_2 & io_storeAddrDone_2; // @[LoadQueue.scala 151:92:@13505.4]
  assign _T_15513 = _T_15512 & addrKnown_15; // @[LoadQueue.scala 152:41:@13506.4]
  assign _T_15514 = addrQ_15 == io_storeAddrQueue_2; // @[LoadQueue.scala 153:30:@13507.4]
  assign conflict_15_2 = _T_15513 & _T_15514; // @[LoadQueue.scala 152:68:@13508.4]
  assign _T_15516 = entriesToCheck_15_3 & io_storeAddrDone_3; // @[LoadQueue.scala 151:92:@13510.4]
  assign _T_15517 = _T_15516 & addrKnown_15; // @[LoadQueue.scala 152:41:@13511.4]
  assign _T_15518 = addrQ_15 == io_storeAddrQueue_3; // @[LoadQueue.scala 153:30:@13512.4]
  assign conflict_15_3 = _T_15517 & _T_15518; // @[LoadQueue.scala 152:68:@13513.4]
  assign _T_15520 = entriesToCheck_15_4 & io_storeAddrDone_4; // @[LoadQueue.scala 151:92:@13515.4]
  assign _T_15521 = _T_15520 & addrKnown_15; // @[LoadQueue.scala 152:41:@13516.4]
  assign _T_15522 = addrQ_15 == io_storeAddrQueue_4; // @[LoadQueue.scala 153:30:@13517.4]
  assign conflict_15_4 = _T_15521 & _T_15522; // @[LoadQueue.scala 152:68:@13518.4]
  assign _T_15524 = entriesToCheck_15_5 & io_storeAddrDone_5; // @[LoadQueue.scala 151:92:@13520.4]
  assign _T_15525 = _T_15524 & addrKnown_15; // @[LoadQueue.scala 152:41:@13521.4]
  assign _T_15526 = addrQ_15 == io_storeAddrQueue_5; // @[LoadQueue.scala 153:30:@13522.4]
  assign conflict_15_5 = _T_15525 & _T_15526; // @[LoadQueue.scala 152:68:@13523.4]
  assign _T_15528 = entriesToCheck_15_6 & io_storeAddrDone_6; // @[LoadQueue.scala 151:92:@13525.4]
  assign _T_15529 = _T_15528 & addrKnown_15; // @[LoadQueue.scala 152:41:@13526.4]
  assign _T_15530 = addrQ_15 == io_storeAddrQueue_6; // @[LoadQueue.scala 153:30:@13527.4]
  assign conflict_15_6 = _T_15529 & _T_15530; // @[LoadQueue.scala 152:68:@13528.4]
  assign _T_15532 = entriesToCheck_15_7 & io_storeAddrDone_7; // @[LoadQueue.scala 151:92:@13530.4]
  assign _T_15533 = _T_15532 & addrKnown_15; // @[LoadQueue.scala 152:41:@13531.4]
  assign _T_15534 = addrQ_15 == io_storeAddrQueue_7; // @[LoadQueue.scala 153:30:@13532.4]
  assign conflict_15_7 = _T_15533 & _T_15534; // @[LoadQueue.scala 152:68:@13533.4]
  assign _T_15536 = entriesToCheck_15_8 & io_storeAddrDone_8; // @[LoadQueue.scala 151:92:@13535.4]
  assign _T_15537 = _T_15536 & addrKnown_15; // @[LoadQueue.scala 152:41:@13536.4]
  assign _T_15538 = addrQ_15 == io_storeAddrQueue_8; // @[LoadQueue.scala 153:30:@13537.4]
  assign conflict_15_8 = _T_15537 & _T_15538; // @[LoadQueue.scala 152:68:@13538.4]
  assign _T_15540 = entriesToCheck_15_9 & io_storeAddrDone_9; // @[LoadQueue.scala 151:92:@13540.4]
  assign _T_15541 = _T_15540 & addrKnown_15; // @[LoadQueue.scala 152:41:@13541.4]
  assign _T_15542 = addrQ_15 == io_storeAddrQueue_9; // @[LoadQueue.scala 153:30:@13542.4]
  assign conflict_15_9 = _T_15541 & _T_15542; // @[LoadQueue.scala 152:68:@13543.4]
  assign _T_15544 = entriesToCheck_15_10 & io_storeAddrDone_10; // @[LoadQueue.scala 151:92:@13545.4]
  assign _T_15545 = _T_15544 & addrKnown_15; // @[LoadQueue.scala 152:41:@13546.4]
  assign _T_15546 = addrQ_15 == io_storeAddrQueue_10; // @[LoadQueue.scala 153:30:@13547.4]
  assign conflict_15_10 = _T_15545 & _T_15546; // @[LoadQueue.scala 152:68:@13548.4]
  assign _T_15548 = entriesToCheck_15_11 & io_storeAddrDone_11; // @[LoadQueue.scala 151:92:@13550.4]
  assign _T_15549 = _T_15548 & addrKnown_15; // @[LoadQueue.scala 152:41:@13551.4]
  assign _T_15550 = addrQ_15 == io_storeAddrQueue_11; // @[LoadQueue.scala 153:30:@13552.4]
  assign conflict_15_11 = _T_15549 & _T_15550; // @[LoadQueue.scala 152:68:@13553.4]
  assign _T_15552 = entriesToCheck_15_12 & io_storeAddrDone_12; // @[LoadQueue.scala 151:92:@13555.4]
  assign _T_15553 = _T_15552 & addrKnown_15; // @[LoadQueue.scala 152:41:@13556.4]
  assign _T_15554 = addrQ_15 == io_storeAddrQueue_12; // @[LoadQueue.scala 153:30:@13557.4]
  assign conflict_15_12 = _T_15553 & _T_15554; // @[LoadQueue.scala 152:68:@13558.4]
  assign _T_15556 = entriesToCheck_15_13 & io_storeAddrDone_13; // @[LoadQueue.scala 151:92:@13560.4]
  assign _T_15557 = _T_15556 & addrKnown_15; // @[LoadQueue.scala 152:41:@13561.4]
  assign _T_15558 = addrQ_15 == io_storeAddrQueue_13; // @[LoadQueue.scala 153:30:@13562.4]
  assign conflict_15_13 = _T_15557 & _T_15558; // @[LoadQueue.scala 152:68:@13563.4]
  assign _T_15560 = entriesToCheck_15_14 & io_storeAddrDone_14; // @[LoadQueue.scala 151:92:@13565.4]
  assign _T_15561 = _T_15560 & addrKnown_15; // @[LoadQueue.scala 152:41:@13566.4]
  assign _T_15562 = addrQ_15 == io_storeAddrQueue_14; // @[LoadQueue.scala 153:30:@13567.4]
  assign conflict_15_14 = _T_15561 & _T_15562; // @[LoadQueue.scala 152:68:@13568.4]
  assign _T_15564 = entriesToCheck_15_15 & io_storeAddrDone_15; // @[LoadQueue.scala 151:92:@13570.4]
  assign _T_15565 = _T_15564 & addrKnown_15; // @[LoadQueue.scala 152:41:@13571.4]
  assign _T_15566 = addrQ_15 == io_storeAddrQueue_15; // @[LoadQueue.scala 153:30:@13572.4]
  assign conflict_15_15 = _T_15565 & _T_15566; // @[LoadQueue.scala 152:68:@13573.4]
  assign _T_16799 = io_storeAddrDone_0 == 1'h0; // @[LoadQueue.scala 163:13:@13576.4]
  assign storeAddrNotKnownFlags_0_0 = _T_16799 & entriesToCheck_0_0; // @[LoadQueue.scala 163:19:@13577.4]
  assign _T_16802 = io_storeAddrDone_1 == 1'h0; // @[LoadQueue.scala 163:13:@13578.4]
  assign storeAddrNotKnownFlags_0_1 = _T_16802 & entriesToCheck_0_1; // @[LoadQueue.scala 163:19:@13579.4]
  assign _T_16805 = io_storeAddrDone_2 == 1'h0; // @[LoadQueue.scala 163:13:@13580.4]
  assign storeAddrNotKnownFlags_0_2 = _T_16805 & entriesToCheck_0_2; // @[LoadQueue.scala 163:19:@13581.4]
  assign _T_16808 = io_storeAddrDone_3 == 1'h0; // @[LoadQueue.scala 163:13:@13582.4]
  assign storeAddrNotKnownFlags_0_3 = _T_16808 & entriesToCheck_0_3; // @[LoadQueue.scala 163:19:@13583.4]
  assign _T_16811 = io_storeAddrDone_4 == 1'h0; // @[LoadQueue.scala 163:13:@13584.4]
  assign storeAddrNotKnownFlags_0_4 = _T_16811 & entriesToCheck_0_4; // @[LoadQueue.scala 163:19:@13585.4]
  assign _T_16814 = io_storeAddrDone_5 == 1'h0; // @[LoadQueue.scala 163:13:@13586.4]
  assign storeAddrNotKnownFlags_0_5 = _T_16814 & entriesToCheck_0_5; // @[LoadQueue.scala 163:19:@13587.4]
  assign _T_16817 = io_storeAddrDone_6 == 1'h0; // @[LoadQueue.scala 163:13:@13588.4]
  assign storeAddrNotKnownFlags_0_6 = _T_16817 & entriesToCheck_0_6; // @[LoadQueue.scala 163:19:@13589.4]
  assign _T_16820 = io_storeAddrDone_7 == 1'h0; // @[LoadQueue.scala 163:13:@13590.4]
  assign storeAddrNotKnownFlags_0_7 = _T_16820 & entriesToCheck_0_7; // @[LoadQueue.scala 163:19:@13591.4]
  assign _T_16823 = io_storeAddrDone_8 == 1'h0; // @[LoadQueue.scala 163:13:@13592.4]
  assign storeAddrNotKnownFlags_0_8 = _T_16823 & entriesToCheck_0_8; // @[LoadQueue.scala 163:19:@13593.4]
  assign _T_16826 = io_storeAddrDone_9 == 1'h0; // @[LoadQueue.scala 163:13:@13594.4]
  assign storeAddrNotKnownFlags_0_9 = _T_16826 & entriesToCheck_0_9; // @[LoadQueue.scala 163:19:@13595.4]
  assign _T_16829 = io_storeAddrDone_10 == 1'h0; // @[LoadQueue.scala 163:13:@13596.4]
  assign storeAddrNotKnownFlags_0_10 = _T_16829 & entriesToCheck_0_10; // @[LoadQueue.scala 163:19:@13597.4]
  assign _T_16832 = io_storeAddrDone_11 == 1'h0; // @[LoadQueue.scala 163:13:@13598.4]
  assign storeAddrNotKnownFlags_0_11 = _T_16832 & entriesToCheck_0_11; // @[LoadQueue.scala 163:19:@13599.4]
  assign _T_16835 = io_storeAddrDone_12 == 1'h0; // @[LoadQueue.scala 163:13:@13600.4]
  assign storeAddrNotKnownFlags_0_12 = _T_16835 & entriesToCheck_0_12; // @[LoadQueue.scala 163:19:@13601.4]
  assign _T_16838 = io_storeAddrDone_13 == 1'h0; // @[LoadQueue.scala 163:13:@13602.4]
  assign storeAddrNotKnownFlags_0_13 = _T_16838 & entriesToCheck_0_13; // @[LoadQueue.scala 163:19:@13603.4]
  assign _T_16841 = io_storeAddrDone_14 == 1'h0; // @[LoadQueue.scala 163:13:@13604.4]
  assign storeAddrNotKnownFlags_0_14 = _T_16841 & entriesToCheck_0_14; // @[LoadQueue.scala 163:19:@13605.4]
  assign _T_16844 = io_storeAddrDone_15 == 1'h0; // @[LoadQueue.scala 163:13:@13606.4]
  assign storeAddrNotKnownFlags_0_15 = _T_16844 & entriesToCheck_0_15; // @[LoadQueue.scala 163:19:@13607.4]
  assign storeAddrNotKnownFlags_1_0 = _T_16799 & entriesToCheck_1_0; // @[LoadQueue.scala 163:19:@13625.4]
  assign storeAddrNotKnownFlags_1_1 = _T_16802 & entriesToCheck_1_1; // @[LoadQueue.scala 163:19:@13627.4]
  assign storeAddrNotKnownFlags_1_2 = _T_16805 & entriesToCheck_1_2; // @[LoadQueue.scala 163:19:@13629.4]
  assign storeAddrNotKnownFlags_1_3 = _T_16808 & entriesToCheck_1_3; // @[LoadQueue.scala 163:19:@13631.4]
  assign storeAddrNotKnownFlags_1_4 = _T_16811 & entriesToCheck_1_4; // @[LoadQueue.scala 163:19:@13633.4]
  assign storeAddrNotKnownFlags_1_5 = _T_16814 & entriesToCheck_1_5; // @[LoadQueue.scala 163:19:@13635.4]
  assign storeAddrNotKnownFlags_1_6 = _T_16817 & entriesToCheck_1_6; // @[LoadQueue.scala 163:19:@13637.4]
  assign storeAddrNotKnownFlags_1_7 = _T_16820 & entriesToCheck_1_7; // @[LoadQueue.scala 163:19:@13639.4]
  assign storeAddrNotKnownFlags_1_8 = _T_16823 & entriesToCheck_1_8; // @[LoadQueue.scala 163:19:@13641.4]
  assign storeAddrNotKnownFlags_1_9 = _T_16826 & entriesToCheck_1_9; // @[LoadQueue.scala 163:19:@13643.4]
  assign storeAddrNotKnownFlags_1_10 = _T_16829 & entriesToCheck_1_10; // @[LoadQueue.scala 163:19:@13645.4]
  assign storeAddrNotKnownFlags_1_11 = _T_16832 & entriesToCheck_1_11; // @[LoadQueue.scala 163:19:@13647.4]
  assign storeAddrNotKnownFlags_1_12 = _T_16835 & entriesToCheck_1_12; // @[LoadQueue.scala 163:19:@13649.4]
  assign storeAddrNotKnownFlags_1_13 = _T_16838 & entriesToCheck_1_13; // @[LoadQueue.scala 163:19:@13651.4]
  assign storeAddrNotKnownFlags_1_14 = _T_16841 & entriesToCheck_1_14; // @[LoadQueue.scala 163:19:@13653.4]
  assign storeAddrNotKnownFlags_1_15 = _T_16844 & entriesToCheck_1_15; // @[LoadQueue.scala 163:19:@13655.4]
  assign storeAddrNotKnownFlags_2_0 = _T_16799 & entriesToCheck_2_0; // @[LoadQueue.scala 163:19:@13673.4]
  assign storeAddrNotKnownFlags_2_1 = _T_16802 & entriesToCheck_2_1; // @[LoadQueue.scala 163:19:@13675.4]
  assign storeAddrNotKnownFlags_2_2 = _T_16805 & entriesToCheck_2_2; // @[LoadQueue.scala 163:19:@13677.4]
  assign storeAddrNotKnownFlags_2_3 = _T_16808 & entriesToCheck_2_3; // @[LoadQueue.scala 163:19:@13679.4]
  assign storeAddrNotKnownFlags_2_4 = _T_16811 & entriesToCheck_2_4; // @[LoadQueue.scala 163:19:@13681.4]
  assign storeAddrNotKnownFlags_2_5 = _T_16814 & entriesToCheck_2_5; // @[LoadQueue.scala 163:19:@13683.4]
  assign storeAddrNotKnownFlags_2_6 = _T_16817 & entriesToCheck_2_6; // @[LoadQueue.scala 163:19:@13685.4]
  assign storeAddrNotKnownFlags_2_7 = _T_16820 & entriesToCheck_2_7; // @[LoadQueue.scala 163:19:@13687.4]
  assign storeAddrNotKnownFlags_2_8 = _T_16823 & entriesToCheck_2_8; // @[LoadQueue.scala 163:19:@13689.4]
  assign storeAddrNotKnownFlags_2_9 = _T_16826 & entriesToCheck_2_9; // @[LoadQueue.scala 163:19:@13691.4]
  assign storeAddrNotKnownFlags_2_10 = _T_16829 & entriesToCheck_2_10; // @[LoadQueue.scala 163:19:@13693.4]
  assign storeAddrNotKnownFlags_2_11 = _T_16832 & entriesToCheck_2_11; // @[LoadQueue.scala 163:19:@13695.4]
  assign storeAddrNotKnownFlags_2_12 = _T_16835 & entriesToCheck_2_12; // @[LoadQueue.scala 163:19:@13697.4]
  assign storeAddrNotKnownFlags_2_13 = _T_16838 & entriesToCheck_2_13; // @[LoadQueue.scala 163:19:@13699.4]
  assign storeAddrNotKnownFlags_2_14 = _T_16841 & entriesToCheck_2_14; // @[LoadQueue.scala 163:19:@13701.4]
  assign storeAddrNotKnownFlags_2_15 = _T_16844 & entriesToCheck_2_15; // @[LoadQueue.scala 163:19:@13703.4]
  assign storeAddrNotKnownFlags_3_0 = _T_16799 & entriesToCheck_3_0; // @[LoadQueue.scala 163:19:@13721.4]
  assign storeAddrNotKnownFlags_3_1 = _T_16802 & entriesToCheck_3_1; // @[LoadQueue.scala 163:19:@13723.4]
  assign storeAddrNotKnownFlags_3_2 = _T_16805 & entriesToCheck_3_2; // @[LoadQueue.scala 163:19:@13725.4]
  assign storeAddrNotKnownFlags_3_3 = _T_16808 & entriesToCheck_3_3; // @[LoadQueue.scala 163:19:@13727.4]
  assign storeAddrNotKnownFlags_3_4 = _T_16811 & entriesToCheck_3_4; // @[LoadQueue.scala 163:19:@13729.4]
  assign storeAddrNotKnownFlags_3_5 = _T_16814 & entriesToCheck_3_5; // @[LoadQueue.scala 163:19:@13731.4]
  assign storeAddrNotKnownFlags_3_6 = _T_16817 & entriesToCheck_3_6; // @[LoadQueue.scala 163:19:@13733.4]
  assign storeAddrNotKnownFlags_3_7 = _T_16820 & entriesToCheck_3_7; // @[LoadQueue.scala 163:19:@13735.4]
  assign storeAddrNotKnownFlags_3_8 = _T_16823 & entriesToCheck_3_8; // @[LoadQueue.scala 163:19:@13737.4]
  assign storeAddrNotKnownFlags_3_9 = _T_16826 & entriesToCheck_3_9; // @[LoadQueue.scala 163:19:@13739.4]
  assign storeAddrNotKnownFlags_3_10 = _T_16829 & entriesToCheck_3_10; // @[LoadQueue.scala 163:19:@13741.4]
  assign storeAddrNotKnownFlags_3_11 = _T_16832 & entriesToCheck_3_11; // @[LoadQueue.scala 163:19:@13743.4]
  assign storeAddrNotKnownFlags_3_12 = _T_16835 & entriesToCheck_3_12; // @[LoadQueue.scala 163:19:@13745.4]
  assign storeAddrNotKnownFlags_3_13 = _T_16838 & entriesToCheck_3_13; // @[LoadQueue.scala 163:19:@13747.4]
  assign storeAddrNotKnownFlags_3_14 = _T_16841 & entriesToCheck_3_14; // @[LoadQueue.scala 163:19:@13749.4]
  assign storeAddrNotKnownFlags_3_15 = _T_16844 & entriesToCheck_3_15; // @[LoadQueue.scala 163:19:@13751.4]
  assign storeAddrNotKnownFlags_4_0 = _T_16799 & entriesToCheck_4_0; // @[LoadQueue.scala 163:19:@13769.4]
  assign storeAddrNotKnownFlags_4_1 = _T_16802 & entriesToCheck_4_1; // @[LoadQueue.scala 163:19:@13771.4]
  assign storeAddrNotKnownFlags_4_2 = _T_16805 & entriesToCheck_4_2; // @[LoadQueue.scala 163:19:@13773.4]
  assign storeAddrNotKnownFlags_4_3 = _T_16808 & entriesToCheck_4_3; // @[LoadQueue.scala 163:19:@13775.4]
  assign storeAddrNotKnownFlags_4_4 = _T_16811 & entriesToCheck_4_4; // @[LoadQueue.scala 163:19:@13777.4]
  assign storeAddrNotKnownFlags_4_5 = _T_16814 & entriesToCheck_4_5; // @[LoadQueue.scala 163:19:@13779.4]
  assign storeAddrNotKnownFlags_4_6 = _T_16817 & entriesToCheck_4_6; // @[LoadQueue.scala 163:19:@13781.4]
  assign storeAddrNotKnownFlags_4_7 = _T_16820 & entriesToCheck_4_7; // @[LoadQueue.scala 163:19:@13783.4]
  assign storeAddrNotKnownFlags_4_8 = _T_16823 & entriesToCheck_4_8; // @[LoadQueue.scala 163:19:@13785.4]
  assign storeAddrNotKnownFlags_4_9 = _T_16826 & entriesToCheck_4_9; // @[LoadQueue.scala 163:19:@13787.4]
  assign storeAddrNotKnownFlags_4_10 = _T_16829 & entriesToCheck_4_10; // @[LoadQueue.scala 163:19:@13789.4]
  assign storeAddrNotKnownFlags_4_11 = _T_16832 & entriesToCheck_4_11; // @[LoadQueue.scala 163:19:@13791.4]
  assign storeAddrNotKnownFlags_4_12 = _T_16835 & entriesToCheck_4_12; // @[LoadQueue.scala 163:19:@13793.4]
  assign storeAddrNotKnownFlags_4_13 = _T_16838 & entriesToCheck_4_13; // @[LoadQueue.scala 163:19:@13795.4]
  assign storeAddrNotKnownFlags_4_14 = _T_16841 & entriesToCheck_4_14; // @[LoadQueue.scala 163:19:@13797.4]
  assign storeAddrNotKnownFlags_4_15 = _T_16844 & entriesToCheck_4_15; // @[LoadQueue.scala 163:19:@13799.4]
  assign storeAddrNotKnownFlags_5_0 = _T_16799 & entriesToCheck_5_0; // @[LoadQueue.scala 163:19:@13817.4]
  assign storeAddrNotKnownFlags_5_1 = _T_16802 & entriesToCheck_5_1; // @[LoadQueue.scala 163:19:@13819.4]
  assign storeAddrNotKnownFlags_5_2 = _T_16805 & entriesToCheck_5_2; // @[LoadQueue.scala 163:19:@13821.4]
  assign storeAddrNotKnownFlags_5_3 = _T_16808 & entriesToCheck_5_3; // @[LoadQueue.scala 163:19:@13823.4]
  assign storeAddrNotKnownFlags_5_4 = _T_16811 & entriesToCheck_5_4; // @[LoadQueue.scala 163:19:@13825.4]
  assign storeAddrNotKnownFlags_5_5 = _T_16814 & entriesToCheck_5_5; // @[LoadQueue.scala 163:19:@13827.4]
  assign storeAddrNotKnownFlags_5_6 = _T_16817 & entriesToCheck_5_6; // @[LoadQueue.scala 163:19:@13829.4]
  assign storeAddrNotKnownFlags_5_7 = _T_16820 & entriesToCheck_5_7; // @[LoadQueue.scala 163:19:@13831.4]
  assign storeAddrNotKnownFlags_5_8 = _T_16823 & entriesToCheck_5_8; // @[LoadQueue.scala 163:19:@13833.4]
  assign storeAddrNotKnownFlags_5_9 = _T_16826 & entriesToCheck_5_9; // @[LoadQueue.scala 163:19:@13835.4]
  assign storeAddrNotKnownFlags_5_10 = _T_16829 & entriesToCheck_5_10; // @[LoadQueue.scala 163:19:@13837.4]
  assign storeAddrNotKnownFlags_5_11 = _T_16832 & entriesToCheck_5_11; // @[LoadQueue.scala 163:19:@13839.4]
  assign storeAddrNotKnownFlags_5_12 = _T_16835 & entriesToCheck_5_12; // @[LoadQueue.scala 163:19:@13841.4]
  assign storeAddrNotKnownFlags_5_13 = _T_16838 & entriesToCheck_5_13; // @[LoadQueue.scala 163:19:@13843.4]
  assign storeAddrNotKnownFlags_5_14 = _T_16841 & entriesToCheck_5_14; // @[LoadQueue.scala 163:19:@13845.4]
  assign storeAddrNotKnownFlags_5_15 = _T_16844 & entriesToCheck_5_15; // @[LoadQueue.scala 163:19:@13847.4]
  assign storeAddrNotKnownFlags_6_0 = _T_16799 & entriesToCheck_6_0; // @[LoadQueue.scala 163:19:@13865.4]
  assign storeAddrNotKnownFlags_6_1 = _T_16802 & entriesToCheck_6_1; // @[LoadQueue.scala 163:19:@13867.4]
  assign storeAddrNotKnownFlags_6_2 = _T_16805 & entriesToCheck_6_2; // @[LoadQueue.scala 163:19:@13869.4]
  assign storeAddrNotKnownFlags_6_3 = _T_16808 & entriesToCheck_6_3; // @[LoadQueue.scala 163:19:@13871.4]
  assign storeAddrNotKnownFlags_6_4 = _T_16811 & entriesToCheck_6_4; // @[LoadQueue.scala 163:19:@13873.4]
  assign storeAddrNotKnownFlags_6_5 = _T_16814 & entriesToCheck_6_5; // @[LoadQueue.scala 163:19:@13875.4]
  assign storeAddrNotKnownFlags_6_6 = _T_16817 & entriesToCheck_6_6; // @[LoadQueue.scala 163:19:@13877.4]
  assign storeAddrNotKnownFlags_6_7 = _T_16820 & entriesToCheck_6_7; // @[LoadQueue.scala 163:19:@13879.4]
  assign storeAddrNotKnownFlags_6_8 = _T_16823 & entriesToCheck_6_8; // @[LoadQueue.scala 163:19:@13881.4]
  assign storeAddrNotKnownFlags_6_9 = _T_16826 & entriesToCheck_6_9; // @[LoadQueue.scala 163:19:@13883.4]
  assign storeAddrNotKnownFlags_6_10 = _T_16829 & entriesToCheck_6_10; // @[LoadQueue.scala 163:19:@13885.4]
  assign storeAddrNotKnownFlags_6_11 = _T_16832 & entriesToCheck_6_11; // @[LoadQueue.scala 163:19:@13887.4]
  assign storeAddrNotKnownFlags_6_12 = _T_16835 & entriesToCheck_6_12; // @[LoadQueue.scala 163:19:@13889.4]
  assign storeAddrNotKnownFlags_6_13 = _T_16838 & entriesToCheck_6_13; // @[LoadQueue.scala 163:19:@13891.4]
  assign storeAddrNotKnownFlags_6_14 = _T_16841 & entriesToCheck_6_14; // @[LoadQueue.scala 163:19:@13893.4]
  assign storeAddrNotKnownFlags_6_15 = _T_16844 & entriesToCheck_6_15; // @[LoadQueue.scala 163:19:@13895.4]
  assign storeAddrNotKnownFlags_7_0 = _T_16799 & entriesToCheck_7_0; // @[LoadQueue.scala 163:19:@13913.4]
  assign storeAddrNotKnownFlags_7_1 = _T_16802 & entriesToCheck_7_1; // @[LoadQueue.scala 163:19:@13915.4]
  assign storeAddrNotKnownFlags_7_2 = _T_16805 & entriesToCheck_7_2; // @[LoadQueue.scala 163:19:@13917.4]
  assign storeAddrNotKnownFlags_7_3 = _T_16808 & entriesToCheck_7_3; // @[LoadQueue.scala 163:19:@13919.4]
  assign storeAddrNotKnownFlags_7_4 = _T_16811 & entriesToCheck_7_4; // @[LoadQueue.scala 163:19:@13921.4]
  assign storeAddrNotKnownFlags_7_5 = _T_16814 & entriesToCheck_7_5; // @[LoadQueue.scala 163:19:@13923.4]
  assign storeAddrNotKnownFlags_7_6 = _T_16817 & entriesToCheck_7_6; // @[LoadQueue.scala 163:19:@13925.4]
  assign storeAddrNotKnownFlags_7_7 = _T_16820 & entriesToCheck_7_7; // @[LoadQueue.scala 163:19:@13927.4]
  assign storeAddrNotKnownFlags_7_8 = _T_16823 & entriesToCheck_7_8; // @[LoadQueue.scala 163:19:@13929.4]
  assign storeAddrNotKnownFlags_7_9 = _T_16826 & entriesToCheck_7_9; // @[LoadQueue.scala 163:19:@13931.4]
  assign storeAddrNotKnownFlags_7_10 = _T_16829 & entriesToCheck_7_10; // @[LoadQueue.scala 163:19:@13933.4]
  assign storeAddrNotKnownFlags_7_11 = _T_16832 & entriesToCheck_7_11; // @[LoadQueue.scala 163:19:@13935.4]
  assign storeAddrNotKnownFlags_7_12 = _T_16835 & entriesToCheck_7_12; // @[LoadQueue.scala 163:19:@13937.4]
  assign storeAddrNotKnownFlags_7_13 = _T_16838 & entriesToCheck_7_13; // @[LoadQueue.scala 163:19:@13939.4]
  assign storeAddrNotKnownFlags_7_14 = _T_16841 & entriesToCheck_7_14; // @[LoadQueue.scala 163:19:@13941.4]
  assign storeAddrNotKnownFlags_7_15 = _T_16844 & entriesToCheck_7_15; // @[LoadQueue.scala 163:19:@13943.4]
  assign storeAddrNotKnownFlags_8_0 = _T_16799 & entriesToCheck_8_0; // @[LoadQueue.scala 163:19:@13961.4]
  assign storeAddrNotKnownFlags_8_1 = _T_16802 & entriesToCheck_8_1; // @[LoadQueue.scala 163:19:@13963.4]
  assign storeAddrNotKnownFlags_8_2 = _T_16805 & entriesToCheck_8_2; // @[LoadQueue.scala 163:19:@13965.4]
  assign storeAddrNotKnownFlags_8_3 = _T_16808 & entriesToCheck_8_3; // @[LoadQueue.scala 163:19:@13967.4]
  assign storeAddrNotKnownFlags_8_4 = _T_16811 & entriesToCheck_8_4; // @[LoadQueue.scala 163:19:@13969.4]
  assign storeAddrNotKnownFlags_8_5 = _T_16814 & entriesToCheck_8_5; // @[LoadQueue.scala 163:19:@13971.4]
  assign storeAddrNotKnownFlags_8_6 = _T_16817 & entriesToCheck_8_6; // @[LoadQueue.scala 163:19:@13973.4]
  assign storeAddrNotKnownFlags_8_7 = _T_16820 & entriesToCheck_8_7; // @[LoadQueue.scala 163:19:@13975.4]
  assign storeAddrNotKnownFlags_8_8 = _T_16823 & entriesToCheck_8_8; // @[LoadQueue.scala 163:19:@13977.4]
  assign storeAddrNotKnownFlags_8_9 = _T_16826 & entriesToCheck_8_9; // @[LoadQueue.scala 163:19:@13979.4]
  assign storeAddrNotKnownFlags_8_10 = _T_16829 & entriesToCheck_8_10; // @[LoadQueue.scala 163:19:@13981.4]
  assign storeAddrNotKnownFlags_8_11 = _T_16832 & entriesToCheck_8_11; // @[LoadQueue.scala 163:19:@13983.4]
  assign storeAddrNotKnownFlags_8_12 = _T_16835 & entriesToCheck_8_12; // @[LoadQueue.scala 163:19:@13985.4]
  assign storeAddrNotKnownFlags_8_13 = _T_16838 & entriesToCheck_8_13; // @[LoadQueue.scala 163:19:@13987.4]
  assign storeAddrNotKnownFlags_8_14 = _T_16841 & entriesToCheck_8_14; // @[LoadQueue.scala 163:19:@13989.4]
  assign storeAddrNotKnownFlags_8_15 = _T_16844 & entriesToCheck_8_15; // @[LoadQueue.scala 163:19:@13991.4]
  assign storeAddrNotKnownFlags_9_0 = _T_16799 & entriesToCheck_9_0; // @[LoadQueue.scala 163:19:@14009.4]
  assign storeAddrNotKnownFlags_9_1 = _T_16802 & entriesToCheck_9_1; // @[LoadQueue.scala 163:19:@14011.4]
  assign storeAddrNotKnownFlags_9_2 = _T_16805 & entriesToCheck_9_2; // @[LoadQueue.scala 163:19:@14013.4]
  assign storeAddrNotKnownFlags_9_3 = _T_16808 & entriesToCheck_9_3; // @[LoadQueue.scala 163:19:@14015.4]
  assign storeAddrNotKnownFlags_9_4 = _T_16811 & entriesToCheck_9_4; // @[LoadQueue.scala 163:19:@14017.4]
  assign storeAddrNotKnownFlags_9_5 = _T_16814 & entriesToCheck_9_5; // @[LoadQueue.scala 163:19:@14019.4]
  assign storeAddrNotKnownFlags_9_6 = _T_16817 & entriesToCheck_9_6; // @[LoadQueue.scala 163:19:@14021.4]
  assign storeAddrNotKnownFlags_9_7 = _T_16820 & entriesToCheck_9_7; // @[LoadQueue.scala 163:19:@14023.4]
  assign storeAddrNotKnownFlags_9_8 = _T_16823 & entriesToCheck_9_8; // @[LoadQueue.scala 163:19:@14025.4]
  assign storeAddrNotKnownFlags_9_9 = _T_16826 & entriesToCheck_9_9; // @[LoadQueue.scala 163:19:@14027.4]
  assign storeAddrNotKnownFlags_9_10 = _T_16829 & entriesToCheck_9_10; // @[LoadQueue.scala 163:19:@14029.4]
  assign storeAddrNotKnownFlags_9_11 = _T_16832 & entriesToCheck_9_11; // @[LoadQueue.scala 163:19:@14031.4]
  assign storeAddrNotKnownFlags_9_12 = _T_16835 & entriesToCheck_9_12; // @[LoadQueue.scala 163:19:@14033.4]
  assign storeAddrNotKnownFlags_9_13 = _T_16838 & entriesToCheck_9_13; // @[LoadQueue.scala 163:19:@14035.4]
  assign storeAddrNotKnownFlags_9_14 = _T_16841 & entriesToCheck_9_14; // @[LoadQueue.scala 163:19:@14037.4]
  assign storeAddrNotKnownFlags_9_15 = _T_16844 & entriesToCheck_9_15; // @[LoadQueue.scala 163:19:@14039.4]
  assign storeAddrNotKnownFlags_10_0 = _T_16799 & entriesToCheck_10_0; // @[LoadQueue.scala 163:19:@14057.4]
  assign storeAddrNotKnownFlags_10_1 = _T_16802 & entriesToCheck_10_1; // @[LoadQueue.scala 163:19:@14059.4]
  assign storeAddrNotKnownFlags_10_2 = _T_16805 & entriesToCheck_10_2; // @[LoadQueue.scala 163:19:@14061.4]
  assign storeAddrNotKnownFlags_10_3 = _T_16808 & entriesToCheck_10_3; // @[LoadQueue.scala 163:19:@14063.4]
  assign storeAddrNotKnownFlags_10_4 = _T_16811 & entriesToCheck_10_4; // @[LoadQueue.scala 163:19:@14065.4]
  assign storeAddrNotKnownFlags_10_5 = _T_16814 & entriesToCheck_10_5; // @[LoadQueue.scala 163:19:@14067.4]
  assign storeAddrNotKnownFlags_10_6 = _T_16817 & entriesToCheck_10_6; // @[LoadQueue.scala 163:19:@14069.4]
  assign storeAddrNotKnownFlags_10_7 = _T_16820 & entriesToCheck_10_7; // @[LoadQueue.scala 163:19:@14071.4]
  assign storeAddrNotKnownFlags_10_8 = _T_16823 & entriesToCheck_10_8; // @[LoadQueue.scala 163:19:@14073.4]
  assign storeAddrNotKnownFlags_10_9 = _T_16826 & entriesToCheck_10_9; // @[LoadQueue.scala 163:19:@14075.4]
  assign storeAddrNotKnownFlags_10_10 = _T_16829 & entriesToCheck_10_10; // @[LoadQueue.scala 163:19:@14077.4]
  assign storeAddrNotKnownFlags_10_11 = _T_16832 & entriesToCheck_10_11; // @[LoadQueue.scala 163:19:@14079.4]
  assign storeAddrNotKnownFlags_10_12 = _T_16835 & entriesToCheck_10_12; // @[LoadQueue.scala 163:19:@14081.4]
  assign storeAddrNotKnownFlags_10_13 = _T_16838 & entriesToCheck_10_13; // @[LoadQueue.scala 163:19:@14083.4]
  assign storeAddrNotKnownFlags_10_14 = _T_16841 & entriesToCheck_10_14; // @[LoadQueue.scala 163:19:@14085.4]
  assign storeAddrNotKnownFlags_10_15 = _T_16844 & entriesToCheck_10_15; // @[LoadQueue.scala 163:19:@14087.4]
  assign storeAddrNotKnownFlags_11_0 = _T_16799 & entriesToCheck_11_0; // @[LoadQueue.scala 163:19:@14105.4]
  assign storeAddrNotKnownFlags_11_1 = _T_16802 & entriesToCheck_11_1; // @[LoadQueue.scala 163:19:@14107.4]
  assign storeAddrNotKnownFlags_11_2 = _T_16805 & entriesToCheck_11_2; // @[LoadQueue.scala 163:19:@14109.4]
  assign storeAddrNotKnownFlags_11_3 = _T_16808 & entriesToCheck_11_3; // @[LoadQueue.scala 163:19:@14111.4]
  assign storeAddrNotKnownFlags_11_4 = _T_16811 & entriesToCheck_11_4; // @[LoadQueue.scala 163:19:@14113.4]
  assign storeAddrNotKnownFlags_11_5 = _T_16814 & entriesToCheck_11_5; // @[LoadQueue.scala 163:19:@14115.4]
  assign storeAddrNotKnownFlags_11_6 = _T_16817 & entriesToCheck_11_6; // @[LoadQueue.scala 163:19:@14117.4]
  assign storeAddrNotKnownFlags_11_7 = _T_16820 & entriesToCheck_11_7; // @[LoadQueue.scala 163:19:@14119.4]
  assign storeAddrNotKnownFlags_11_8 = _T_16823 & entriesToCheck_11_8; // @[LoadQueue.scala 163:19:@14121.4]
  assign storeAddrNotKnownFlags_11_9 = _T_16826 & entriesToCheck_11_9; // @[LoadQueue.scala 163:19:@14123.4]
  assign storeAddrNotKnownFlags_11_10 = _T_16829 & entriesToCheck_11_10; // @[LoadQueue.scala 163:19:@14125.4]
  assign storeAddrNotKnownFlags_11_11 = _T_16832 & entriesToCheck_11_11; // @[LoadQueue.scala 163:19:@14127.4]
  assign storeAddrNotKnownFlags_11_12 = _T_16835 & entriesToCheck_11_12; // @[LoadQueue.scala 163:19:@14129.4]
  assign storeAddrNotKnownFlags_11_13 = _T_16838 & entriesToCheck_11_13; // @[LoadQueue.scala 163:19:@14131.4]
  assign storeAddrNotKnownFlags_11_14 = _T_16841 & entriesToCheck_11_14; // @[LoadQueue.scala 163:19:@14133.4]
  assign storeAddrNotKnownFlags_11_15 = _T_16844 & entriesToCheck_11_15; // @[LoadQueue.scala 163:19:@14135.4]
  assign storeAddrNotKnownFlags_12_0 = _T_16799 & entriesToCheck_12_0; // @[LoadQueue.scala 163:19:@14153.4]
  assign storeAddrNotKnownFlags_12_1 = _T_16802 & entriesToCheck_12_1; // @[LoadQueue.scala 163:19:@14155.4]
  assign storeAddrNotKnownFlags_12_2 = _T_16805 & entriesToCheck_12_2; // @[LoadQueue.scala 163:19:@14157.4]
  assign storeAddrNotKnownFlags_12_3 = _T_16808 & entriesToCheck_12_3; // @[LoadQueue.scala 163:19:@14159.4]
  assign storeAddrNotKnownFlags_12_4 = _T_16811 & entriesToCheck_12_4; // @[LoadQueue.scala 163:19:@14161.4]
  assign storeAddrNotKnownFlags_12_5 = _T_16814 & entriesToCheck_12_5; // @[LoadQueue.scala 163:19:@14163.4]
  assign storeAddrNotKnownFlags_12_6 = _T_16817 & entriesToCheck_12_6; // @[LoadQueue.scala 163:19:@14165.4]
  assign storeAddrNotKnownFlags_12_7 = _T_16820 & entriesToCheck_12_7; // @[LoadQueue.scala 163:19:@14167.4]
  assign storeAddrNotKnownFlags_12_8 = _T_16823 & entriesToCheck_12_8; // @[LoadQueue.scala 163:19:@14169.4]
  assign storeAddrNotKnownFlags_12_9 = _T_16826 & entriesToCheck_12_9; // @[LoadQueue.scala 163:19:@14171.4]
  assign storeAddrNotKnownFlags_12_10 = _T_16829 & entriesToCheck_12_10; // @[LoadQueue.scala 163:19:@14173.4]
  assign storeAddrNotKnownFlags_12_11 = _T_16832 & entriesToCheck_12_11; // @[LoadQueue.scala 163:19:@14175.4]
  assign storeAddrNotKnownFlags_12_12 = _T_16835 & entriesToCheck_12_12; // @[LoadQueue.scala 163:19:@14177.4]
  assign storeAddrNotKnownFlags_12_13 = _T_16838 & entriesToCheck_12_13; // @[LoadQueue.scala 163:19:@14179.4]
  assign storeAddrNotKnownFlags_12_14 = _T_16841 & entriesToCheck_12_14; // @[LoadQueue.scala 163:19:@14181.4]
  assign storeAddrNotKnownFlags_12_15 = _T_16844 & entriesToCheck_12_15; // @[LoadQueue.scala 163:19:@14183.4]
  assign storeAddrNotKnownFlags_13_0 = _T_16799 & entriesToCheck_13_0; // @[LoadQueue.scala 163:19:@14201.4]
  assign storeAddrNotKnownFlags_13_1 = _T_16802 & entriesToCheck_13_1; // @[LoadQueue.scala 163:19:@14203.4]
  assign storeAddrNotKnownFlags_13_2 = _T_16805 & entriesToCheck_13_2; // @[LoadQueue.scala 163:19:@14205.4]
  assign storeAddrNotKnownFlags_13_3 = _T_16808 & entriesToCheck_13_3; // @[LoadQueue.scala 163:19:@14207.4]
  assign storeAddrNotKnownFlags_13_4 = _T_16811 & entriesToCheck_13_4; // @[LoadQueue.scala 163:19:@14209.4]
  assign storeAddrNotKnownFlags_13_5 = _T_16814 & entriesToCheck_13_5; // @[LoadQueue.scala 163:19:@14211.4]
  assign storeAddrNotKnownFlags_13_6 = _T_16817 & entriesToCheck_13_6; // @[LoadQueue.scala 163:19:@14213.4]
  assign storeAddrNotKnownFlags_13_7 = _T_16820 & entriesToCheck_13_7; // @[LoadQueue.scala 163:19:@14215.4]
  assign storeAddrNotKnownFlags_13_8 = _T_16823 & entriesToCheck_13_8; // @[LoadQueue.scala 163:19:@14217.4]
  assign storeAddrNotKnownFlags_13_9 = _T_16826 & entriesToCheck_13_9; // @[LoadQueue.scala 163:19:@14219.4]
  assign storeAddrNotKnownFlags_13_10 = _T_16829 & entriesToCheck_13_10; // @[LoadQueue.scala 163:19:@14221.4]
  assign storeAddrNotKnownFlags_13_11 = _T_16832 & entriesToCheck_13_11; // @[LoadQueue.scala 163:19:@14223.4]
  assign storeAddrNotKnownFlags_13_12 = _T_16835 & entriesToCheck_13_12; // @[LoadQueue.scala 163:19:@14225.4]
  assign storeAddrNotKnownFlags_13_13 = _T_16838 & entriesToCheck_13_13; // @[LoadQueue.scala 163:19:@14227.4]
  assign storeAddrNotKnownFlags_13_14 = _T_16841 & entriesToCheck_13_14; // @[LoadQueue.scala 163:19:@14229.4]
  assign storeAddrNotKnownFlags_13_15 = _T_16844 & entriesToCheck_13_15; // @[LoadQueue.scala 163:19:@14231.4]
  assign storeAddrNotKnownFlags_14_0 = _T_16799 & entriesToCheck_14_0; // @[LoadQueue.scala 163:19:@14249.4]
  assign storeAddrNotKnownFlags_14_1 = _T_16802 & entriesToCheck_14_1; // @[LoadQueue.scala 163:19:@14251.4]
  assign storeAddrNotKnownFlags_14_2 = _T_16805 & entriesToCheck_14_2; // @[LoadQueue.scala 163:19:@14253.4]
  assign storeAddrNotKnownFlags_14_3 = _T_16808 & entriesToCheck_14_3; // @[LoadQueue.scala 163:19:@14255.4]
  assign storeAddrNotKnownFlags_14_4 = _T_16811 & entriesToCheck_14_4; // @[LoadQueue.scala 163:19:@14257.4]
  assign storeAddrNotKnownFlags_14_5 = _T_16814 & entriesToCheck_14_5; // @[LoadQueue.scala 163:19:@14259.4]
  assign storeAddrNotKnownFlags_14_6 = _T_16817 & entriesToCheck_14_6; // @[LoadQueue.scala 163:19:@14261.4]
  assign storeAddrNotKnownFlags_14_7 = _T_16820 & entriesToCheck_14_7; // @[LoadQueue.scala 163:19:@14263.4]
  assign storeAddrNotKnownFlags_14_8 = _T_16823 & entriesToCheck_14_8; // @[LoadQueue.scala 163:19:@14265.4]
  assign storeAddrNotKnownFlags_14_9 = _T_16826 & entriesToCheck_14_9; // @[LoadQueue.scala 163:19:@14267.4]
  assign storeAddrNotKnownFlags_14_10 = _T_16829 & entriesToCheck_14_10; // @[LoadQueue.scala 163:19:@14269.4]
  assign storeAddrNotKnownFlags_14_11 = _T_16832 & entriesToCheck_14_11; // @[LoadQueue.scala 163:19:@14271.4]
  assign storeAddrNotKnownFlags_14_12 = _T_16835 & entriesToCheck_14_12; // @[LoadQueue.scala 163:19:@14273.4]
  assign storeAddrNotKnownFlags_14_13 = _T_16838 & entriesToCheck_14_13; // @[LoadQueue.scala 163:19:@14275.4]
  assign storeAddrNotKnownFlags_14_14 = _T_16841 & entriesToCheck_14_14; // @[LoadQueue.scala 163:19:@14277.4]
  assign storeAddrNotKnownFlags_14_15 = _T_16844 & entriesToCheck_14_15; // @[LoadQueue.scala 163:19:@14279.4]
  assign storeAddrNotKnownFlags_15_0 = _T_16799 & entriesToCheck_15_0; // @[LoadQueue.scala 163:19:@14297.4]
  assign storeAddrNotKnownFlags_15_1 = _T_16802 & entriesToCheck_15_1; // @[LoadQueue.scala 163:19:@14299.4]
  assign storeAddrNotKnownFlags_15_2 = _T_16805 & entriesToCheck_15_2; // @[LoadQueue.scala 163:19:@14301.4]
  assign storeAddrNotKnownFlags_15_3 = _T_16808 & entriesToCheck_15_3; // @[LoadQueue.scala 163:19:@14303.4]
  assign storeAddrNotKnownFlags_15_4 = _T_16811 & entriesToCheck_15_4; // @[LoadQueue.scala 163:19:@14305.4]
  assign storeAddrNotKnownFlags_15_5 = _T_16814 & entriesToCheck_15_5; // @[LoadQueue.scala 163:19:@14307.4]
  assign storeAddrNotKnownFlags_15_6 = _T_16817 & entriesToCheck_15_6; // @[LoadQueue.scala 163:19:@14309.4]
  assign storeAddrNotKnownFlags_15_7 = _T_16820 & entriesToCheck_15_7; // @[LoadQueue.scala 163:19:@14311.4]
  assign storeAddrNotKnownFlags_15_8 = _T_16823 & entriesToCheck_15_8; // @[LoadQueue.scala 163:19:@14313.4]
  assign storeAddrNotKnownFlags_15_9 = _T_16826 & entriesToCheck_15_9; // @[LoadQueue.scala 163:19:@14315.4]
  assign storeAddrNotKnownFlags_15_10 = _T_16829 & entriesToCheck_15_10; // @[LoadQueue.scala 163:19:@14317.4]
  assign storeAddrNotKnownFlags_15_11 = _T_16832 & entriesToCheck_15_11; // @[LoadQueue.scala 163:19:@14319.4]
  assign storeAddrNotKnownFlags_15_12 = _T_16835 & entriesToCheck_15_12; // @[LoadQueue.scala 163:19:@14321.4]
  assign storeAddrNotKnownFlags_15_13 = _T_16838 & entriesToCheck_15_13; // @[LoadQueue.scala 163:19:@14323.4]
  assign storeAddrNotKnownFlags_15_14 = _T_16841 & entriesToCheck_15_14; // @[LoadQueue.scala 163:19:@14325.4]
  assign storeAddrNotKnownFlags_15_15 = _T_16844 & entriesToCheck_15_15; // @[LoadQueue.scala 163:19:@14327.4]
  assign _T_18002 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@14658.4]
  assign _T_18009 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8}; // @[Mux.scala 19:72:@14665.4]
  assign _T_18010 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,_T_18002}; // @[Mux.scala 19:72:@14666.4]
  assign _T_18012 = _T_2689 ? _T_18010 : 16'h0; // @[Mux.scala 19:72:@14667.4]
  assign _T_18019 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@14674.4]
  assign _T_18026 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9}; // @[Mux.scala 19:72:@14681.4]
  assign _T_18027 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,_T_18019}; // @[Mux.scala 19:72:@14682.4]
  assign _T_18029 = _T_2690 ? _T_18027 : 16'h0; // @[Mux.scala 19:72:@14683.4]
  assign _T_18036 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@14690.4]
  assign _T_18043 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10}; // @[Mux.scala 19:72:@14697.4]
  assign _T_18044 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,_T_18036}; // @[Mux.scala 19:72:@14698.4]
  assign _T_18046 = _T_2691 ? _T_18044 : 16'h0; // @[Mux.scala 19:72:@14699.4]
  assign _T_18053 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@14706.4]
  assign _T_18060 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11}; // @[Mux.scala 19:72:@14713.4]
  assign _T_18061 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,_T_18053}; // @[Mux.scala 19:72:@14714.4]
  assign _T_18063 = _T_2692 ? _T_18061 : 16'h0; // @[Mux.scala 19:72:@14715.4]
  assign _T_18070 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@14722.4]
  assign _T_18077 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12}; // @[Mux.scala 19:72:@14729.4]
  assign _T_18078 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,_T_18070}; // @[Mux.scala 19:72:@14730.4]
  assign _T_18080 = _T_2693 ? _T_18078 : 16'h0; // @[Mux.scala 19:72:@14731.4]
  assign _T_18087 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@14738.4]
  assign _T_18094 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13}; // @[Mux.scala 19:72:@14745.4]
  assign _T_18095 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,_T_18087}; // @[Mux.scala 19:72:@14746.4]
  assign _T_18097 = _T_2694 ? _T_18095 : 16'h0; // @[Mux.scala 19:72:@14747.4]
  assign _T_18104 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@14754.4]
  assign _T_18111 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14}; // @[Mux.scala 19:72:@14761.4]
  assign _T_18112 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,_T_18104}; // @[Mux.scala 19:72:@14762.4]
  assign _T_18114 = _T_2695 ? _T_18112 : 16'h0; // @[Mux.scala 19:72:@14763.4]
  assign _T_18121 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7}; // @[Mux.scala 19:72:@14770.4]
  assign _T_18128 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15}; // @[Mux.scala 19:72:@14777.4]
  assign _T_18129 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,_T_18121}; // @[Mux.scala 19:72:@14778.4]
  assign _T_18131 = _T_2696 ? _T_18129 : 16'h0; // @[Mux.scala 19:72:@14779.4]
  assign _T_18146 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,_T_18009}; // @[Mux.scala 19:72:@14794.4]
  assign _T_18148 = _T_2697 ? _T_18146 : 16'h0; // @[Mux.scala 19:72:@14795.4]
  assign _T_18163 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,_T_18026}; // @[Mux.scala 19:72:@14810.4]
  assign _T_18165 = _T_2698 ? _T_18163 : 16'h0; // @[Mux.scala 19:72:@14811.4]
  assign _T_18180 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,_T_18043}; // @[Mux.scala 19:72:@14826.4]
  assign _T_18182 = _T_2699 ? _T_18180 : 16'h0; // @[Mux.scala 19:72:@14827.4]
  assign _T_18197 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,_T_18060}; // @[Mux.scala 19:72:@14842.4]
  assign _T_18199 = _T_2700 ? _T_18197 : 16'h0; // @[Mux.scala 19:72:@14843.4]
  assign _T_18214 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,_T_18077}; // @[Mux.scala 19:72:@14858.4]
  assign _T_18216 = _T_2701 ? _T_18214 : 16'h0; // @[Mux.scala 19:72:@14859.4]
  assign _T_18231 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,_T_18094}; // @[Mux.scala 19:72:@14874.4]
  assign _T_18233 = _T_2702 ? _T_18231 : 16'h0; // @[Mux.scala 19:72:@14875.4]
  assign _T_18248 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,_T_18111}; // @[Mux.scala 19:72:@14890.4]
  assign _T_18250 = _T_2703 ? _T_18248 : 16'h0; // @[Mux.scala 19:72:@14891.4]
  assign _T_18265 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,_T_18128}; // @[Mux.scala 19:72:@14906.4]
  assign _T_18267 = _T_2704 ? _T_18265 : 16'h0; // @[Mux.scala 19:72:@14907.4]
  assign _T_18268 = _T_18012 | _T_18029; // @[Mux.scala 19:72:@14908.4]
  assign _T_18269 = _T_18268 | _T_18046; // @[Mux.scala 19:72:@14909.4]
  assign _T_18270 = _T_18269 | _T_18063; // @[Mux.scala 19:72:@14910.4]
  assign _T_18271 = _T_18270 | _T_18080; // @[Mux.scala 19:72:@14911.4]
  assign _T_18272 = _T_18271 | _T_18097; // @[Mux.scala 19:72:@14912.4]
  assign _T_18273 = _T_18272 | _T_18114; // @[Mux.scala 19:72:@14913.4]
  assign _T_18274 = _T_18273 | _T_18131; // @[Mux.scala 19:72:@14914.4]
  assign _T_18275 = _T_18274 | _T_18148; // @[Mux.scala 19:72:@14915.4]
  assign _T_18276 = _T_18275 | _T_18165; // @[Mux.scala 19:72:@14916.4]
  assign _T_18277 = _T_18276 | _T_18182; // @[Mux.scala 19:72:@14917.4]
  assign _T_18278 = _T_18277 | _T_18199; // @[Mux.scala 19:72:@14918.4]
  assign _T_18279 = _T_18278 | _T_18216; // @[Mux.scala 19:72:@14919.4]
  assign _T_18280 = _T_18279 | _T_18233; // @[Mux.scala 19:72:@14920.4]
  assign _T_18281 = _T_18280 | _T_18250; // @[Mux.scala 19:72:@14921.4]
  assign _T_18282 = _T_18281 | _T_18267; // @[Mux.scala 19:72:@14922.4]
  assign _T_18860 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@15272.4]
  assign _T_18867 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8}; // @[Mux.scala 19:72:@15279.4]
  assign _T_18868 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,_T_18860}; // @[Mux.scala 19:72:@15280.4]
  assign _T_18870 = _T_2689 ? _T_18868 : 16'h0; // @[Mux.scala 19:72:@15281.4]
  assign _T_18877 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@15288.4]
  assign _T_18884 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9}; // @[Mux.scala 19:72:@15295.4]
  assign _T_18885 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,_T_18877}; // @[Mux.scala 19:72:@15296.4]
  assign _T_18887 = _T_2690 ? _T_18885 : 16'h0; // @[Mux.scala 19:72:@15297.4]
  assign _T_18894 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@15304.4]
  assign _T_18901 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10}; // @[Mux.scala 19:72:@15311.4]
  assign _T_18902 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,_T_18894}; // @[Mux.scala 19:72:@15312.4]
  assign _T_18904 = _T_2691 ? _T_18902 : 16'h0; // @[Mux.scala 19:72:@15313.4]
  assign _T_18911 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@15320.4]
  assign _T_18918 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11}; // @[Mux.scala 19:72:@15327.4]
  assign _T_18919 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,_T_18911}; // @[Mux.scala 19:72:@15328.4]
  assign _T_18921 = _T_2692 ? _T_18919 : 16'h0; // @[Mux.scala 19:72:@15329.4]
  assign _T_18928 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@15336.4]
  assign _T_18935 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12}; // @[Mux.scala 19:72:@15343.4]
  assign _T_18936 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,_T_18928}; // @[Mux.scala 19:72:@15344.4]
  assign _T_18938 = _T_2693 ? _T_18936 : 16'h0; // @[Mux.scala 19:72:@15345.4]
  assign _T_18945 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@15352.4]
  assign _T_18952 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13}; // @[Mux.scala 19:72:@15359.4]
  assign _T_18953 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,_T_18945}; // @[Mux.scala 19:72:@15360.4]
  assign _T_18955 = _T_2694 ? _T_18953 : 16'h0; // @[Mux.scala 19:72:@15361.4]
  assign _T_18962 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@15368.4]
  assign _T_18969 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14}; // @[Mux.scala 19:72:@15375.4]
  assign _T_18970 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,_T_18962}; // @[Mux.scala 19:72:@15376.4]
  assign _T_18972 = _T_2695 ? _T_18970 : 16'h0; // @[Mux.scala 19:72:@15377.4]
  assign _T_18979 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7}; // @[Mux.scala 19:72:@15384.4]
  assign _T_18986 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15}; // @[Mux.scala 19:72:@15391.4]
  assign _T_18987 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,_T_18979}; // @[Mux.scala 19:72:@15392.4]
  assign _T_18989 = _T_2696 ? _T_18987 : 16'h0; // @[Mux.scala 19:72:@15393.4]
  assign _T_19004 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,_T_18867}; // @[Mux.scala 19:72:@15408.4]
  assign _T_19006 = _T_2697 ? _T_19004 : 16'h0; // @[Mux.scala 19:72:@15409.4]
  assign _T_19021 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,_T_18884}; // @[Mux.scala 19:72:@15424.4]
  assign _T_19023 = _T_2698 ? _T_19021 : 16'h0; // @[Mux.scala 19:72:@15425.4]
  assign _T_19038 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,_T_18901}; // @[Mux.scala 19:72:@15440.4]
  assign _T_19040 = _T_2699 ? _T_19038 : 16'h0; // @[Mux.scala 19:72:@15441.4]
  assign _T_19055 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,_T_18918}; // @[Mux.scala 19:72:@15456.4]
  assign _T_19057 = _T_2700 ? _T_19055 : 16'h0; // @[Mux.scala 19:72:@15457.4]
  assign _T_19072 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,_T_18935}; // @[Mux.scala 19:72:@15472.4]
  assign _T_19074 = _T_2701 ? _T_19072 : 16'h0; // @[Mux.scala 19:72:@15473.4]
  assign _T_19089 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,_T_18952}; // @[Mux.scala 19:72:@15488.4]
  assign _T_19091 = _T_2702 ? _T_19089 : 16'h0; // @[Mux.scala 19:72:@15489.4]
  assign _T_19106 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,_T_18969}; // @[Mux.scala 19:72:@15504.4]
  assign _T_19108 = _T_2703 ? _T_19106 : 16'h0; // @[Mux.scala 19:72:@15505.4]
  assign _T_19123 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,_T_18986}; // @[Mux.scala 19:72:@15520.4]
  assign _T_19125 = _T_2704 ? _T_19123 : 16'h0; // @[Mux.scala 19:72:@15521.4]
  assign _T_19126 = _T_18870 | _T_18887; // @[Mux.scala 19:72:@15522.4]
  assign _T_19127 = _T_19126 | _T_18904; // @[Mux.scala 19:72:@15523.4]
  assign _T_19128 = _T_19127 | _T_18921; // @[Mux.scala 19:72:@15524.4]
  assign _T_19129 = _T_19128 | _T_18938; // @[Mux.scala 19:72:@15525.4]
  assign _T_19130 = _T_19129 | _T_18955; // @[Mux.scala 19:72:@15526.4]
  assign _T_19131 = _T_19130 | _T_18972; // @[Mux.scala 19:72:@15527.4]
  assign _T_19132 = _T_19131 | _T_18989; // @[Mux.scala 19:72:@15528.4]
  assign _T_19133 = _T_19132 | _T_19006; // @[Mux.scala 19:72:@15529.4]
  assign _T_19134 = _T_19133 | _T_19023; // @[Mux.scala 19:72:@15530.4]
  assign _T_19135 = _T_19134 | _T_19040; // @[Mux.scala 19:72:@15531.4]
  assign _T_19136 = _T_19135 | _T_19057; // @[Mux.scala 19:72:@15532.4]
  assign _T_19137 = _T_19136 | _T_19074; // @[Mux.scala 19:72:@15533.4]
  assign _T_19138 = _T_19137 | _T_19091; // @[Mux.scala 19:72:@15534.4]
  assign _T_19139 = _T_19138 | _T_19108; // @[Mux.scala 19:72:@15535.4]
  assign _T_19140 = _T_19139 | _T_19125; // @[Mux.scala 19:72:@15536.4]
  assign _T_19718 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@15886.4]
  assign _T_19725 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8}; // @[Mux.scala 19:72:@15893.4]
  assign _T_19726 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,_T_19718}; // @[Mux.scala 19:72:@15894.4]
  assign _T_19728 = _T_2689 ? _T_19726 : 16'h0; // @[Mux.scala 19:72:@15895.4]
  assign _T_19735 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@15902.4]
  assign _T_19742 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9}; // @[Mux.scala 19:72:@15909.4]
  assign _T_19743 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,_T_19735}; // @[Mux.scala 19:72:@15910.4]
  assign _T_19745 = _T_2690 ? _T_19743 : 16'h0; // @[Mux.scala 19:72:@15911.4]
  assign _T_19752 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@15918.4]
  assign _T_19759 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10}; // @[Mux.scala 19:72:@15925.4]
  assign _T_19760 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,_T_19752}; // @[Mux.scala 19:72:@15926.4]
  assign _T_19762 = _T_2691 ? _T_19760 : 16'h0; // @[Mux.scala 19:72:@15927.4]
  assign _T_19769 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@15934.4]
  assign _T_19776 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11}; // @[Mux.scala 19:72:@15941.4]
  assign _T_19777 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,_T_19769}; // @[Mux.scala 19:72:@15942.4]
  assign _T_19779 = _T_2692 ? _T_19777 : 16'h0; // @[Mux.scala 19:72:@15943.4]
  assign _T_19786 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@15950.4]
  assign _T_19793 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12}; // @[Mux.scala 19:72:@15957.4]
  assign _T_19794 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,_T_19786}; // @[Mux.scala 19:72:@15958.4]
  assign _T_19796 = _T_2693 ? _T_19794 : 16'h0; // @[Mux.scala 19:72:@15959.4]
  assign _T_19803 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@15966.4]
  assign _T_19810 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13}; // @[Mux.scala 19:72:@15973.4]
  assign _T_19811 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,_T_19803}; // @[Mux.scala 19:72:@15974.4]
  assign _T_19813 = _T_2694 ? _T_19811 : 16'h0; // @[Mux.scala 19:72:@15975.4]
  assign _T_19820 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@15982.4]
  assign _T_19827 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14}; // @[Mux.scala 19:72:@15989.4]
  assign _T_19828 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,_T_19820}; // @[Mux.scala 19:72:@15990.4]
  assign _T_19830 = _T_2695 ? _T_19828 : 16'h0; // @[Mux.scala 19:72:@15991.4]
  assign _T_19837 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7}; // @[Mux.scala 19:72:@15998.4]
  assign _T_19844 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15}; // @[Mux.scala 19:72:@16005.4]
  assign _T_19845 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,_T_19837}; // @[Mux.scala 19:72:@16006.4]
  assign _T_19847 = _T_2696 ? _T_19845 : 16'h0; // @[Mux.scala 19:72:@16007.4]
  assign _T_19862 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,_T_19725}; // @[Mux.scala 19:72:@16022.4]
  assign _T_19864 = _T_2697 ? _T_19862 : 16'h0; // @[Mux.scala 19:72:@16023.4]
  assign _T_19879 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,_T_19742}; // @[Mux.scala 19:72:@16038.4]
  assign _T_19881 = _T_2698 ? _T_19879 : 16'h0; // @[Mux.scala 19:72:@16039.4]
  assign _T_19896 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,_T_19759}; // @[Mux.scala 19:72:@16054.4]
  assign _T_19898 = _T_2699 ? _T_19896 : 16'h0; // @[Mux.scala 19:72:@16055.4]
  assign _T_19913 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,_T_19776}; // @[Mux.scala 19:72:@16070.4]
  assign _T_19915 = _T_2700 ? _T_19913 : 16'h0; // @[Mux.scala 19:72:@16071.4]
  assign _T_19930 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,_T_19793}; // @[Mux.scala 19:72:@16086.4]
  assign _T_19932 = _T_2701 ? _T_19930 : 16'h0; // @[Mux.scala 19:72:@16087.4]
  assign _T_19947 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,_T_19810}; // @[Mux.scala 19:72:@16102.4]
  assign _T_19949 = _T_2702 ? _T_19947 : 16'h0; // @[Mux.scala 19:72:@16103.4]
  assign _T_19964 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,_T_19827}; // @[Mux.scala 19:72:@16118.4]
  assign _T_19966 = _T_2703 ? _T_19964 : 16'h0; // @[Mux.scala 19:72:@16119.4]
  assign _T_19981 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,_T_19844}; // @[Mux.scala 19:72:@16134.4]
  assign _T_19983 = _T_2704 ? _T_19981 : 16'h0; // @[Mux.scala 19:72:@16135.4]
  assign _T_19984 = _T_19728 | _T_19745; // @[Mux.scala 19:72:@16136.4]
  assign _T_19985 = _T_19984 | _T_19762; // @[Mux.scala 19:72:@16137.4]
  assign _T_19986 = _T_19985 | _T_19779; // @[Mux.scala 19:72:@16138.4]
  assign _T_19987 = _T_19986 | _T_19796; // @[Mux.scala 19:72:@16139.4]
  assign _T_19988 = _T_19987 | _T_19813; // @[Mux.scala 19:72:@16140.4]
  assign _T_19989 = _T_19988 | _T_19830; // @[Mux.scala 19:72:@16141.4]
  assign _T_19990 = _T_19989 | _T_19847; // @[Mux.scala 19:72:@16142.4]
  assign _T_19991 = _T_19990 | _T_19864; // @[Mux.scala 19:72:@16143.4]
  assign _T_19992 = _T_19991 | _T_19881; // @[Mux.scala 19:72:@16144.4]
  assign _T_19993 = _T_19992 | _T_19898; // @[Mux.scala 19:72:@16145.4]
  assign _T_19994 = _T_19993 | _T_19915; // @[Mux.scala 19:72:@16146.4]
  assign _T_19995 = _T_19994 | _T_19932; // @[Mux.scala 19:72:@16147.4]
  assign _T_19996 = _T_19995 | _T_19949; // @[Mux.scala 19:72:@16148.4]
  assign _T_19997 = _T_19996 | _T_19966; // @[Mux.scala 19:72:@16149.4]
  assign _T_19998 = _T_19997 | _T_19983; // @[Mux.scala 19:72:@16150.4]
  assign _T_20576 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@16500.4]
  assign _T_20583 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8}; // @[Mux.scala 19:72:@16507.4]
  assign _T_20584 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,_T_20576}; // @[Mux.scala 19:72:@16508.4]
  assign _T_20586 = _T_2689 ? _T_20584 : 16'h0; // @[Mux.scala 19:72:@16509.4]
  assign _T_20593 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@16516.4]
  assign _T_20600 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9}; // @[Mux.scala 19:72:@16523.4]
  assign _T_20601 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,_T_20593}; // @[Mux.scala 19:72:@16524.4]
  assign _T_20603 = _T_2690 ? _T_20601 : 16'h0; // @[Mux.scala 19:72:@16525.4]
  assign _T_20610 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@16532.4]
  assign _T_20617 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10}; // @[Mux.scala 19:72:@16539.4]
  assign _T_20618 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,_T_20610}; // @[Mux.scala 19:72:@16540.4]
  assign _T_20620 = _T_2691 ? _T_20618 : 16'h0; // @[Mux.scala 19:72:@16541.4]
  assign _T_20627 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@16548.4]
  assign _T_20634 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11}; // @[Mux.scala 19:72:@16555.4]
  assign _T_20635 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,_T_20627}; // @[Mux.scala 19:72:@16556.4]
  assign _T_20637 = _T_2692 ? _T_20635 : 16'h0; // @[Mux.scala 19:72:@16557.4]
  assign _T_20644 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@16564.4]
  assign _T_20651 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12}; // @[Mux.scala 19:72:@16571.4]
  assign _T_20652 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,_T_20644}; // @[Mux.scala 19:72:@16572.4]
  assign _T_20654 = _T_2693 ? _T_20652 : 16'h0; // @[Mux.scala 19:72:@16573.4]
  assign _T_20661 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@16580.4]
  assign _T_20668 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13}; // @[Mux.scala 19:72:@16587.4]
  assign _T_20669 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,_T_20661}; // @[Mux.scala 19:72:@16588.4]
  assign _T_20671 = _T_2694 ? _T_20669 : 16'h0; // @[Mux.scala 19:72:@16589.4]
  assign _T_20678 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@16596.4]
  assign _T_20685 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14}; // @[Mux.scala 19:72:@16603.4]
  assign _T_20686 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,_T_20678}; // @[Mux.scala 19:72:@16604.4]
  assign _T_20688 = _T_2695 ? _T_20686 : 16'h0; // @[Mux.scala 19:72:@16605.4]
  assign _T_20695 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7}; // @[Mux.scala 19:72:@16612.4]
  assign _T_20702 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15}; // @[Mux.scala 19:72:@16619.4]
  assign _T_20703 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,_T_20695}; // @[Mux.scala 19:72:@16620.4]
  assign _T_20705 = _T_2696 ? _T_20703 : 16'h0; // @[Mux.scala 19:72:@16621.4]
  assign _T_20720 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,_T_20583}; // @[Mux.scala 19:72:@16636.4]
  assign _T_20722 = _T_2697 ? _T_20720 : 16'h0; // @[Mux.scala 19:72:@16637.4]
  assign _T_20737 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,_T_20600}; // @[Mux.scala 19:72:@16652.4]
  assign _T_20739 = _T_2698 ? _T_20737 : 16'h0; // @[Mux.scala 19:72:@16653.4]
  assign _T_20754 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,_T_20617}; // @[Mux.scala 19:72:@16668.4]
  assign _T_20756 = _T_2699 ? _T_20754 : 16'h0; // @[Mux.scala 19:72:@16669.4]
  assign _T_20771 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,_T_20634}; // @[Mux.scala 19:72:@16684.4]
  assign _T_20773 = _T_2700 ? _T_20771 : 16'h0; // @[Mux.scala 19:72:@16685.4]
  assign _T_20788 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,_T_20651}; // @[Mux.scala 19:72:@16700.4]
  assign _T_20790 = _T_2701 ? _T_20788 : 16'h0; // @[Mux.scala 19:72:@16701.4]
  assign _T_20805 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,_T_20668}; // @[Mux.scala 19:72:@16716.4]
  assign _T_20807 = _T_2702 ? _T_20805 : 16'h0; // @[Mux.scala 19:72:@16717.4]
  assign _T_20822 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,_T_20685}; // @[Mux.scala 19:72:@16732.4]
  assign _T_20824 = _T_2703 ? _T_20822 : 16'h0; // @[Mux.scala 19:72:@16733.4]
  assign _T_20839 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,_T_20702}; // @[Mux.scala 19:72:@16748.4]
  assign _T_20841 = _T_2704 ? _T_20839 : 16'h0; // @[Mux.scala 19:72:@16749.4]
  assign _T_20842 = _T_20586 | _T_20603; // @[Mux.scala 19:72:@16750.4]
  assign _T_20843 = _T_20842 | _T_20620; // @[Mux.scala 19:72:@16751.4]
  assign _T_20844 = _T_20843 | _T_20637; // @[Mux.scala 19:72:@16752.4]
  assign _T_20845 = _T_20844 | _T_20654; // @[Mux.scala 19:72:@16753.4]
  assign _T_20846 = _T_20845 | _T_20671; // @[Mux.scala 19:72:@16754.4]
  assign _T_20847 = _T_20846 | _T_20688; // @[Mux.scala 19:72:@16755.4]
  assign _T_20848 = _T_20847 | _T_20705; // @[Mux.scala 19:72:@16756.4]
  assign _T_20849 = _T_20848 | _T_20722; // @[Mux.scala 19:72:@16757.4]
  assign _T_20850 = _T_20849 | _T_20739; // @[Mux.scala 19:72:@16758.4]
  assign _T_20851 = _T_20850 | _T_20756; // @[Mux.scala 19:72:@16759.4]
  assign _T_20852 = _T_20851 | _T_20773; // @[Mux.scala 19:72:@16760.4]
  assign _T_20853 = _T_20852 | _T_20790; // @[Mux.scala 19:72:@16761.4]
  assign _T_20854 = _T_20853 | _T_20807; // @[Mux.scala 19:72:@16762.4]
  assign _T_20855 = _T_20854 | _T_20824; // @[Mux.scala 19:72:@16763.4]
  assign _T_20856 = _T_20855 | _T_20841; // @[Mux.scala 19:72:@16764.4]
  assign _T_21434 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@17114.4]
  assign _T_21441 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8}; // @[Mux.scala 19:72:@17121.4]
  assign _T_21442 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,_T_21434}; // @[Mux.scala 19:72:@17122.4]
  assign _T_21444 = _T_2689 ? _T_21442 : 16'h0; // @[Mux.scala 19:72:@17123.4]
  assign _T_21451 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@17130.4]
  assign _T_21458 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9}; // @[Mux.scala 19:72:@17137.4]
  assign _T_21459 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,_T_21451}; // @[Mux.scala 19:72:@17138.4]
  assign _T_21461 = _T_2690 ? _T_21459 : 16'h0; // @[Mux.scala 19:72:@17139.4]
  assign _T_21468 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@17146.4]
  assign _T_21475 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10}; // @[Mux.scala 19:72:@17153.4]
  assign _T_21476 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,_T_21468}; // @[Mux.scala 19:72:@17154.4]
  assign _T_21478 = _T_2691 ? _T_21476 : 16'h0; // @[Mux.scala 19:72:@17155.4]
  assign _T_21485 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@17162.4]
  assign _T_21492 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11}; // @[Mux.scala 19:72:@17169.4]
  assign _T_21493 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,_T_21485}; // @[Mux.scala 19:72:@17170.4]
  assign _T_21495 = _T_2692 ? _T_21493 : 16'h0; // @[Mux.scala 19:72:@17171.4]
  assign _T_21502 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@17178.4]
  assign _T_21509 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12}; // @[Mux.scala 19:72:@17185.4]
  assign _T_21510 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,_T_21502}; // @[Mux.scala 19:72:@17186.4]
  assign _T_21512 = _T_2693 ? _T_21510 : 16'h0; // @[Mux.scala 19:72:@17187.4]
  assign _T_21519 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@17194.4]
  assign _T_21526 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13}; // @[Mux.scala 19:72:@17201.4]
  assign _T_21527 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,_T_21519}; // @[Mux.scala 19:72:@17202.4]
  assign _T_21529 = _T_2694 ? _T_21527 : 16'h0; // @[Mux.scala 19:72:@17203.4]
  assign _T_21536 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@17210.4]
  assign _T_21543 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14}; // @[Mux.scala 19:72:@17217.4]
  assign _T_21544 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,_T_21536}; // @[Mux.scala 19:72:@17218.4]
  assign _T_21546 = _T_2695 ? _T_21544 : 16'h0; // @[Mux.scala 19:72:@17219.4]
  assign _T_21553 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7}; // @[Mux.scala 19:72:@17226.4]
  assign _T_21560 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15}; // @[Mux.scala 19:72:@17233.4]
  assign _T_21561 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,_T_21553}; // @[Mux.scala 19:72:@17234.4]
  assign _T_21563 = _T_2696 ? _T_21561 : 16'h0; // @[Mux.scala 19:72:@17235.4]
  assign _T_21578 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,_T_21441}; // @[Mux.scala 19:72:@17250.4]
  assign _T_21580 = _T_2697 ? _T_21578 : 16'h0; // @[Mux.scala 19:72:@17251.4]
  assign _T_21595 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,_T_21458}; // @[Mux.scala 19:72:@17266.4]
  assign _T_21597 = _T_2698 ? _T_21595 : 16'h0; // @[Mux.scala 19:72:@17267.4]
  assign _T_21612 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,_T_21475}; // @[Mux.scala 19:72:@17282.4]
  assign _T_21614 = _T_2699 ? _T_21612 : 16'h0; // @[Mux.scala 19:72:@17283.4]
  assign _T_21629 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,_T_21492}; // @[Mux.scala 19:72:@17298.4]
  assign _T_21631 = _T_2700 ? _T_21629 : 16'h0; // @[Mux.scala 19:72:@17299.4]
  assign _T_21646 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,_T_21509}; // @[Mux.scala 19:72:@17314.4]
  assign _T_21648 = _T_2701 ? _T_21646 : 16'h0; // @[Mux.scala 19:72:@17315.4]
  assign _T_21663 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,_T_21526}; // @[Mux.scala 19:72:@17330.4]
  assign _T_21665 = _T_2702 ? _T_21663 : 16'h0; // @[Mux.scala 19:72:@17331.4]
  assign _T_21680 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,_T_21543}; // @[Mux.scala 19:72:@17346.4]
  assign _T_21682 = _T_2703 ? _T_21680 : 16'h0; // @[Mux.scala 19:72:@17347.4]
  assign _T_21697 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,_T_21560}; // @[Mux.scala 19:72:@17362.4]
  assign _T_21699 = _T_2704 ? _T_21697 : 16'h0; // @[Mux.scala 19:72:@17363.4]
  assign _T_21700 = _T_21444 | _T_21461; // @[Mux.scala 19:72:@17364.4]
  assign _T_21701 = _T_21700 | _T_21478; // @[Mux.scala 19:72:@17365.4]
  assign _T_21702 = _T_21701 | _T_21495; // @[Mux.scala 19:72:@17366.4]
  assign _T_21703 = _T_21702 | _T_21512; // @[Mux.scala 19:72:@17367.4]
  assign _T_21704 = _T_21703 | _T_21529; // @[Mux.scala 19:72:@17368.4]
  assign _T_21705 = _T_21704 | _T_21546; // @[Mux.scala 19:72:@17369.4]
  assign _T_21706 = _T_21705 | _T_21563; // @[Mux.scala 19:72:@17370.4]
  assign _T_21707 = _T_21706 | _T_21580; // @[Mux.scala 19:72:@17371.4]
  assign _T_21708 = _T_21707 | _T_21597; // @[Mux.scala 19:72:@17372.4]
  assign _T_21709 = _T_21708 | _T_21614; // @[Mux.scala 19:72:@17373.4]
  assign _T_21710 = _T_21709 | _T_21631; // @[Mux.scala 19:72:@17374.4]
  assign _T_21711 = _T_21710 | _T_21648; // @[Mux.scala 19:72:@17375.4]
  assign _T_21712 = _T_21711 | _T_21665; // @[Mux.scala 19:72:@17376.4]
  assign _T_21713 = _T_21712 | _T_21682; // @[Mux.scala 19:72:@17377.4]
  assign _T_21714 = _T_21713 | _T_21699; // @[Mux.scala 19:72:@17378.4]
  assign _T_22292 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@17728.4]
  assign _T_22299 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8}; // @[Mux.scala 19:72:@17735.4]
  assign _T_22300 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,_T_22292}; // @[Mux.scala 19:72:@17736.4]
  assign _T_22302 = _T_2689 ? _T_22300 : 16'h0; // @[Mux.scala 19:72:@17737.4]
  assign _T_22309 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@17744.4]
  assign _T_22316 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9}; // @[Mux.scala 19:72:@17751.4]
  assign _T_22317 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,_T_22309}; // @[Mux.scala 19:72:@17752.4]
  assign _T_22319 = _T_2690 ? _T_22317 : 16'h0; // @[Mux.scala 19:72:@17753.4]
  assign _T_22326 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@17760.4]
  assign _T_22333 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10}; // @[Mux.scala 19:72:@17767.4]
  assign _T_22334 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,_T_22326}; // @[Mux.scala 19:72:@17768.4]
  assign _T_22336 = _T_2691 ? _T_22334 : 16'h0; // @[Mux.scala 19:72:@17769.4]
  assign _T_22343 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@17776.4]
  assign _T_22350 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11}; // @[Mux.scala 19:72:@17783.4]
  assign _T_22351 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,_T_22343}; // @[Mux.scala 19:72:@17784.4]
  assign _T_22353 = _T_2692 ? _T_22351 : 16'h0; // @[Mux.scala 19:72:@17785.4]
  assign _T_22360 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@17792.4]
  assign _T_22367 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12}; // @[Mux.scala 19:72:@17799.4]
  assign _T_22368 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,_T_22360}; // @[Mux.scala 19:72:@17800.4]
  assign _T_22370 = _T_2693 ? _T_22368 : 16'h0; // @[Mux.scala 19:72:@17801.4]
  assign _T_22377 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@17808.4]
  assign _T_22384 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13}; // @[Mux.scala 19:72:@17815.4]
  assign _T_22385 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,_T_22377}; // @[Mux.scala 19:72:@17816.4]
  assign _T_22387 = _T_2694 ? _T_22385 : 16'h0; // @[Mux.scala 19:72:@17817.4]
  assign _T_22394 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@17824.4]
  assign _T_22401 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14}; // @[Mux.scala 19:72:@17831.4]
  assign _T_22402 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,_T_22394}; // @[Mux.scala 19:72:@17832.4]
  assign _T_22404 = _T_2695 ? _T_22402 : 16'h0; // @[Mux.scala 19:72:@17833.4]
  assign _T_22411 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7}; // @[Mux.scala 19:72:@17840.4]
  assign _T_22418 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15}; // @[Mux.scala 19:72:@17847.4]
  assign _T_22419 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,_T_22411}; // @[Mux.scala 19:72:@17848.4]
  assign _T_22421 = _T_2696 ? _T_22419 : 16'h0; // @[Mux.scala 19:72:@17849.4]
  assign _T_22436 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,_T_22299}; // @[Mux.scala 19:72:@17864.4]
  assign _T_22438 = _T_2697 ? _T_22436 : 16'h0; // @[Mux.scala 19:72:@17865.4]
  assign _T_22453 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,_T_22316}; // @[Mux.scala 19:72:@17880.4]
  assign _T_22455 = _T_2698 ? _T_22453 : 16'h0; // @[Mux.scala 19:72:@17881.4]
  assign _T_22470 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,_T_22333}; // @[Mux.scala 19:72:@17896.4]
  assign _T_22472 = _T_2699 ? _T_22470 : 16'h0; // @[Mux.scala 19:72:@17897.4]
  assign _T_22487 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,_T_22350}; // @[Mux.scala 19:72:@17912.4]
  assign _T_22489 = _T_2700 ? _T_22487 : 16'h0; // @[Mux.scala 19:72:@17913.4]
  assign _T_22504 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,_T_22367}; // @[Mux.scala 19:72:@17928.4]
  assign _T_22506 = _T_2701 ? _T_22504 : 16'h0; // @[Mux.scala 19:72:@17929.4]
  assign _T_22521 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,_T_22384}; // @[Mux.scala 19:72:@17944.4]
  assign _T_22523 = _T_2702 ? _T_22521 : 16'h0; // @[Mux.scala 19:72:@17945.4]
  assign _T_22538 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,_T_22401}; // @[Mux.scala 19:72:@17960.4]
  assign _T_22540 = _T_2703 ? _T_22538 : 16'h0; // @[Mux.scala 19:72:@17961.4]
  assign _T_22555 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,_T_22418}; // @[Mux.scala 19:72:@17976.4]
  assign _T_22557 = _T_2704 ? _T_22555 : 16'h0; // @[Mux.scala 19:72:@17977.4]
  assign _T_22558 = _T_22302 | _T_22319; // @[Mux.scala 19:72:@17978.4]
  assign _T_22559 = _T_22558 | _T_22336; // @[Mux.scala 19:72:@17979.4]
  assign _T_22560 = _T_22559 | _T_22353; // @[Mux.scala 19:72:@17980.4]
  assign _T_22561 = _T_22560 | _T_22370; // @[Mux.scala 19:72:@17981.4]
  assign _T_22562 = _T_22561 | _T_22387; // @[Mux.scala 19:72:@17982.4]
  assign _T_22563 = _T_22562 | _T_22404; // @[Mux.scala 19:72:@17983.4]
  assign _T_22564 = _T_22563 | _T_22421; // @[Mux.scala 19:72:@17984.4]
  assign _T_22565 = _T_22564 | _T_22438; // @[Mux.scala 19:72:@17985.4]
  assign _T_22566 = _T_22565 | _T_22455; // @[Mux.scala 19:72:@17986.4]
  assign _T_22567 = _T_22566 | _T_22472; // @[Mux.scala 19:72:@17987.4]
  assign _T_22568 = _T_22567 | _T_22489; // @[Mux.scala 19:72:@17988.4]
  assign _T_22569 = _T_22568 | _T_22506; // @[Mux.scala 19:72:@17989.4]
  assign _T_22570 = _T_22569 | _T_22523; // @[Mux.scala 19:72:@17990.4]
  assign _T_22571 = _T_22570 | _T_22540; // @[Mux.scala 19:72:@17991.4]
  assign _T_22572 = _T_22571 | _T_22557; // @[Mux.scala 19:72:@17992.4]
  assign _T_23150 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@18342.4]
  assign _T_23157 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8}; // @[Mux.scala 19:72:@18349.4]
  assign _T_23158 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,_T_23150}; // @[Mux.scala 19:72:@18350.4]
  assign _T_23160 = _T_2689 ? _T_23158 : 16'h0; // @[Mux.scala 19:72:@18351.4]
  assign _T_23167 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@18358.4]
  assign _T_23174 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9}; // @[Mux.scala 19:72:@18365.4]
  assign _T_23175 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,_T_23167}; // @[Mux.scala 19:72:@18366.4]
  assign _T_23177 = _T_2690 ? _T_23175 : 16'h0; // @[Mux.scala 19:72:@18367.4]
  assign _T_23184 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@18374.4]
  assign _T_23191 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10}; // @[Mux.scala 19:72:@18381.4]
  assign _T_23192 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,_T_23184}; // @[Mux.scala 19:72:@18382.4]
  assign _T_23194 = _T_2691 ? _T_23192 : 16'h0; // @[Mux.scala 19:72:@18383.4]
  assign _T_23201 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@18390.4]
  assign _T_23208 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11}; // @[Mux.scala 19:72:@18397.4]
  assign _T_23209 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,_T_23201}; // @[Mux.scala 19:72:@18398.4]
  assign _T_23211 = _T_2692 ? _T_23209 : 16'h0; // @[Mux.scala 19:72:@18399.4]
  assign _T_23218 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@18406.4]
  assign _T_23225 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12}; // @[Mux.scala 19:72:@18413.4]
  assign _T_23226 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,_T_23218}; // @[Mux.scala 19:72:@18414.4]
  assign _T_23228 = _T_2693 ? _T_23226 : 16'h0; // @[Mux.scala 19:72:@18415.4]
  assign _T_23235 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@18422.4]
  assign _T_23242 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13}; // @[Mux.scala 19:72:@18429.4]
  assign _T_23243 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,_T_23235}; // @[Mux.scala 19:72:@18430.4]
  assign _T_23245 = _T_2694 ? _T_23243 : 16'h0; // @[Mux.scala 19:72:@18431.4]
  assign _T_23252 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@18438.4]
  assign _T_23259 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14}; // @[Mux.scala 19:72:@18445.4]
  assign _T_23260 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,_T_23252}; // @[Mux.scala 19:72:@18446.4]
  assign _T_23262 = _T_2695 ? _T_23260 : 16'h0; // @[Mux.scala 19:72:@18447.4]
  assign _T_23269 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7}; // @[Mux.scala 19:72:@18454.4]
  assign _T_23276 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15}; // @[Mux.scala 19:72:@18461.4]
  assign _T_23277 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,_T_23269}; // @[Mux.scala 19:72:@18462.4]
  assign _T_23279 = _T_2696 ? _T_23277 : 16'h0; // @[Mux.scala 19:72:@18463.4]
  assign _T_23294 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,_T_23157}; // @[Mux.scala 19:72:@18478.4]
  assign _T_23296 = _T_2697 ? _T_23294 : 16'h0; // @[Mux.scala 19:72:@18479.4]
  assign _T_23311 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,_T_23174}; // @[Mux.scala 19:72:@18494.4]
  assign _T_23313 = _T_2698 ? _T_23311 : 16'h0; // @[Mux.scala 19:72:@18495.4]
  assign _T_23328 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,_T_23191}; // @[Mux.scala 19:72:@18510.4]
  assign _T_23330 = _T_2699 ? _T_23328 : 16'h0; // @[Mux.scala 19:72:@18511.4]
  assign _T_23345 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,_T_23208}; // @[Mux.scala 19:72:@18526.4]
  assign _T_23347 = _T_2700 ? _T_23345 : 16'h0; // @[Mux.scala 19:72:@18527.4]
  assign _T_23362 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,_T_23225}; // @[Mux.scala 19:72:@18542.4]
  assign _T_23364 = _T_2701 ? _T_23362 : 16'h0; // @[Mux.scala 19:72:@18543.4]
  assign _T_23379 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,_T_23242}; // @[Mux.scala 19:72:@18558.4]
  assign _T_23381 = _T_2702 ? _T_23379 : 16'h0; // @[Mux.scala 19:72:@18559.4]
  assign _T_23396 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,_T_23259}; // @[Mux.scala 19:72:@18574.4]
  assign _T_23398 = _T_2703 ? _T_23396 : 16'h0; // @[Mux.scala 19:72:@18575.4]
  assign _T_23413 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,_T_23276}; // @[Mux.scala 19:72:@18590.4]
  assign _T_23415 = _T_2704 ? _T_23413 : 16'h0; // @[Mux.scala 19:72:@18591.4]
  assign _T_23416 = _T_23160 | _T_23177; // @[Mux.scala 19:72:@18592.4]
  assign _T_23417 = _T_23416 | _T_23194; // @[Mux.scala 19:72:@18593.4]
  assign _T_23418 = _T_23417 | _T_23211; // @[Mux.scala 19:72:@18594.4]
  assign _T_23419 = _T_23418 | _T_23228; // @[Mux.scala 19:72:@18595.4]
  assign _T_23420 = _T_23419 | _T_23245; // @[Mux.scala 19:72:@18596.4]
  assign _T_23421 = _T_23420 | _T_23262; // @[Mux.scala 19:72:@18597.4]
  assign _T_23422 = _T_23421 | _T_23279; // @[Mux.scala 19:72:@18598.4]
  assign _T_23423 = _T_23422 | _T_23296; // @[Mux.scala 19:72:@18599.4]
  assign _T_23424 = _T_23423 | _T_23313; // @[Mux.scala 19:72:@18600.4]
  assign _T_23425 = _T_23424 | _T_23330; // @[Mux.scala 19:72:@18601.4]
  assign _T_23426 = _T_23425 | _T_23347; // @[Mux.scala 19:72:@18602.4]
  assign _T_23427 = _T_23426 | _T_23364; // @[Mux.scala 19:72:@18603.4]
  assign _T_23428 = _T_23427 | _T_23381; // @[Mux.scala 19:72:@18604.4]
  assign _T_23429 = _T_23428 | _T_23398; // @[Mux.scala 19:72:@18605.4]
  assign _T_23430 = _T_23429 | _T_23415; // @[Mux.scala 19:72:@18606.4]
  assign _T_24008 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@18956.4]
  assign _T_24015 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8}; // @[Mux.scala 19:72:@18963.4]
  assign _T_24016 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,_T_24008}; // @[Mux.scala 19:72:@18964.4]
  assign _T_24018 = _T_2689 ? _T_24016 : 16'h0; // @[Mux.scala 19:72:@18965.4]
  assign _T_24025 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@18972.4]
  assign _T_24032 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9}; // @[Mux.scala 19:72:@18979.4]
  assign _T_24033 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,_T_24025}; // @[Mux.scala 19:72:@18980.4]
  assign _T_24035 = _T_2690 ? _T_24033 : 16'h0; // @[Mux.scala 19:72:@18981.4]
  assign _T_24042 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@18988.4]
  assign _T_24049 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10}; // @[Mux.scala 19:72:@18995.4]
  assign _T_24050 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,_T_24042}; // @[Mux.scala 19:72:@18996.4]
  assign _T_24052 = _T_2691 ? _T_24050 : 16'h0; // @[Mux.scala 19:72:@18997.4]
  assign _T_24059 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@19004.4]
  assign _T_24066 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11}; // @[Mux.scala 19:72:@19011.4]
  assign _T_24067 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,_T_24059}; // @[Mux.scala 19:72:@19012.4]
  assign _T_24069 = _T_2692 ? _T_24067 : 16'h0; // @[Mux.scala 19:72:@19013.4]
  assign _T_24076 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@19020.4]
  assign _T_24083 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12}; // @[Mux.scala 19:72:@19027.4]
  assign _T_24084 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,_T_24076}; // @[Mux.scala 19:72:@19028.4]
  assign _T_24086 = _T_2693 ? _T_24084 : 16'h0; // @[Mux.scala 19:72:@19029.4]
  assign _T_24093 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@19036.4]
  assign _T_24100 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13}; // @[Mux.scala 19:72:@19043.4]
  assign _T_24101 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,_T_24093}; // @[Mux.scala 19:72:@19044.4]
  assign _T_24103 = _T_2694 ? _T_24101 : 16'h0; // @[Mux.scala 19:72:@19045.4]
  assign _T_24110 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@19052.4]
  assign _T_24117 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14}; // @[Mux.scala 19:72:@19059.4]
  assign _T_24118 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,_T_24110}; // @[Mux.scala 19:72:@19060.4]
  assign _T_24120 = _T_2695 ? _T_24118 : 16'h0; // @[Mux.scala 19:72:@19061.4]
  assign _T_24127 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7}; // @[Mux.scala 19:72:@19068.4]
  assign _T_24134 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15}; // @[Mux.scala 19:72:@19075.4]
  assign _T_24135 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,_T_24127}; // @[Mux.scala 19:72:@19076.4]
  assign _T_24137 = _T_2696 ? _T_24135 : 16'h0; // @[Mux.scala 19:72:@19077.4]
  assign _T_24152 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,_T_24015}; // @[Mux.scala 19:72:@19092.4]
  assign _T_24154 = _T_2697 ? _T_24152 : 16'h0; // @[Mux.scala 19:72:@19093.4]
  assign _T_24169 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,_T_24032}; // @[Mux.scala 19:72:@19108.4]
  assign _T_24171 = _T_2698 ? _T_24169 : 16'h0; // @[Mux.scala 19:72:@19109.4]
  assign _T_24186 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,_T_24049}; // @[Mux.scala 19:72:@19124.4]
  assign _T_24188 = _T_2699 ? _T_24186 : 16'h0; // @[Mux.scala 19:72:@19125.4]
  assign _T_24203 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,_T_24066}; // @[Mux.scala 19:72:@19140.4]
  assign _T_24205 = _T_2700 ? _T_24203 : 16'h0; // @[Mux.scala 19:72:@19141.4]
  assign _T_24220 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,_T_24083}; // @[Mux.scala 19:72:@19156.4]
  assign _T_24222 = _T_2701 ? _T_24220 : 16'h0; // @[Mux.scala 19:72:@19157.4]
  assign _T_24237 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,_T_24100}; // @[Mux.scala 19:72:@19172.4]
  assign _T_24239 = _T_2702 ? _T_24237 : 16'h0; // @[Mux.scala 19:72:@19173.4]
  assign _T_24254 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,_T_24117}; // @[Mux.scala 19:72:@19188.4]
  assign _T_24256 = _T_2703 ? _T_24254 : 16'h0; // @[Mux.scala 19:72:@19189.4]
  assign _T_24271 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,_T_24134}; // @[Mux.scala 19:72:@19204.4]
  assign _T_24273 = _T_2704 ? _T_24271 : 16'h0; // @[Mux.scala 19:72:@19205.4]
  assign _T_24274 = _T_24018 | _T_24035; // @[Mux.scala 19:72:@19206.4]
  assign _T_24275 = _T_24274 | _T_24052; // @[Mux.scala 19:72:@19207.4]
  assign _T_24276 = _T_24275 | _T_24069; // @[Mux.scala 19:72:@19208.4]
  assign _T_24277 = _T_24276 | _T_24086; // @[Mux.scala 19:72:@19209.4]
  assign _T_24278 = _T_24277 | _T_24103; // @[Mux.scala 19:72:@19210.4]
  assign _T_24279 = _T_24278 | _T_24120; // @[Mux.scala 19:72:@19211.4]
  assign _T_24280 = _T_24279 | _T_24137; // @[Mux.scala 19:72:@19212.4]
  assign _T_24281 = _T_24280 | _T_24154; // @[Mux.scala 19:72:@19213.4]
  assign _T_24282 = _T_24281 | _T_24171; // @[Mux.scala 19:72:@19214.4]
  assign _T_24283 = _T_24282 | _T_24188; // @[Mux.scala 19:72:@19215.4]
  assign _T_24284 = _T_24283 | _T_24205; // @[Mux.scala 19:72:@19216.4]
  assign _T_24285 = _T_24284 | _T_24222; // @[Mux.scala 19:72:@19217.4]
  assign _T_24286 = _T_24285 | _T_24239; // @[Mux.scala 19:72:@19218.4]
  assign _T_24287 = _T_24286 | _T_24256; // @[Mux.scala 19:72:@19219.4]
  assign _T_24288 = _T_24287 | _T_24273; // @[Mux.scala 19:72:@19220.4]
  assign _T_24866 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0}; // @[Mux.scala 19:72:@19570.4]
  assign _T_24873 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8}; // @[Mux.scala 19:72:@19577.4]
  assign _T_24874 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,_T_24866}; // @[Mux.scala 19:72:@19578.4]
  assign _T_24876 = _T_2689 ? _T_24874 : 16'h0; // @[Mux.scala 19:72:@19579.4]
  assign _T_24883 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1}; // @[Mux.scala 19:72:@19586.4]
  assign _T_24890 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9}; // @[Mux.scala 19:72:@19593.4]
  assign _T_24891 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,_T_24883}; // @[Mux.scala 19:72:@19594.4]
  assign _T_24893 = _T_2690 ? _T_24891 : 16'h0; // @[Mux.scala 19:72:@19595.4]
  assign _T_24900 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2}; // @[Mux.scala 19:72:@19602.4]
  assign _T_24907 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10}; // @[Mux.scala 19:72:@19609.4]
  assign _T_24908 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,_T_24900}; // @[Mux.scala 19:72:@19610.4]
  assign _T_24910 = _T_2691 ? _T_24908 : 16'h0; // @[Mux.scala 19:72:@19611.4]
  assign _T_24917 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3}; // @[Mux.scala 19:72:@19618.4]
  assign _T_24924 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11}; // @[Mux.scala 19:72:@19625.4]
  assign _T_24925 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,_T_24917}; // @[Mux.scala 19:72:@19626.4]
  assign _T_24927 = _T_2692 ? _T_24925 : 16'h0; // @[Mux.scala 19:72:@19627.4]
  assign _T_24934 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4}; // @[Mux.scala 19:72:@19634.4]
  assign _T_24941 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12}; // @[Mux.scala 19:72:@19641.4]
  assign _T_24942 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,_T_24934}; // @[Mux.scala 19:72:@19642.4]
  assign _T_24944 = _T_2693 ? _T_24942 : 16'h0; // @[Mux.scala 19:72:@19643.4]
  assign _T_24951 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5}; // @[Mux.scala 19:72:@19650.4]
  assign _T_24958 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13}; // @[Mux.scala 19:72:@19657.4]
  assign _T_24959 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,_T_24951}; // @[Mux.scala 19:72:@19658.4]
  assign _T_24961 = _T_2694 ? _T_24959 : 16'h0; // @[Mux.scala 19:72:@19659.4]
  assign _T_24968 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6}; // @[Mux.scala 19:72:@19666.4]
  assign _T_24975 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14}; // @[Mux.scala 19:72:@19673.4]
  assign _T_24976 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,_T_24968}; // @[Mux.scala 19:72:@19674.4]
  assign _T_24978 = _T_2695 ? _T_24976 : 16'h0; // @[Mux.scala 19:72:@19675.4]
  assign _T_24985 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7}; // @[Mux.scala 19:72:@19682.4]
  assign _T_24992 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15}; // @[Mux.scala 19:72:@19689.4]
  assign _T_24993 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,_T_24985}; // @[Mux.scala 19:72:@19690.4]
  assign _T_24995 = _T_2696 ? _T_24993 : 16'h0; // @[Mux.scala 19:72:@19691.4]
  assign _T_25010 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,_T_24873}; // @[Mux.scala 19:72:@19706.4]
  assign _T_25012 = _T_2697 ? _T_25010 : 16'h0; // @[Mux.scala 19:72:@19707.4]
  assign _T_25027 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,_T_24890}; // @[Mux.scala 19:72:@19722.4]
  assign _T_25029 = _T_2698 ? _T_25027 : 16'h0; // @[Mux.scala 19:72:@19723.4]
  assign _T_25044 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,_T_24907}; // @[Mux.scala 19:72:@19738.4]
  assign _T_25046 = _T_2699 ? _T_25044 : 16'h0; // @[Mux.scala 19:72:@19739.4]
  assign _T_25061 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,_T_24924}; // @[Mux.scala 19:72:@19754.4]
  assign _T_25063 = _T_2700 ? _T_25061 : 16'h0; // @[Mux.scala 19:72:@19755.4]
  assign _T_25078 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,_T_24941}; // @[Mux.scala 19:72:@19770.4]
  assign _T_25080 = _T_2701 ? _T_25078 : 16'h0; // @[Mux.scala 19:72:@19771.4]
  assign _T_25095 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,_T_24958}; // @[Mux.scala 19:72:@19786.4]
  assign _T_25097 = _T_2702 ? _T_25095 : 16'h0; // @[Mux.scala 19:72:@19787.4]
  assign _T_25112 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,_T_24975}; // @[Mux.scala 19:72:@19802.4]
  assign _T_25114 = _T_2703 ? _T_25112 : 16'h0; // @[Mux.scala 19:72:@19803.4]
  assign _T_25129 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,_T_24992}; // @[Mux.scala 19:72:@19818.4]
  assign _T_25131 = _T_2704 ? _T_25129 : 16'h0; // @[Mux.scala 19:72:@19819.4]
  assign _T_25132 = _T_24876 | _T_24893; // @[Mux.scala 19:72:@19820.4]
  assign _T_25133 = _T_25132 | _T_24910; // @[Mux.scala 19:72:@19821.4]
  assign _T_25134 = _T_25133 | _T_24927; // @[Mux.scala 19:72:@19822.4]
  assign _T_25135 = _T_25134 | _T_24944; // @[Mux.scala 19:72:@19823.4]
  assign _T_25136 = _T_25135 | _T_24961; // @[Mux.scala 19:72:@19824.4]
  assign _T_25137 = _T_25136 | _T_24978; // @[Mux.scala 19:72:@19825.4]
  assign _T_25138 = _T_25137 | _T_24995; // @[Mux.scala 19:72:@19826.4]
  assign _T_25139 = _T_25138 | _T_25012; // @[Mux.scala 19:72:@19827.4]
  assign _T_25140 = _T_25139 | _T_25029; // @[Mux.scala 19:72:@19828.4]
  assign _T_25141 = _T_25140 | _T_25046; // @[Mux.scala 19:72:@19829.4]
  assign _T_25142 = _T_25141 | _T_25063; // @[Mux.scala 19:72:@19830.4]
  assign _T_25143 = _T_25142 | _T_25080; // @[Mux.scala 19:72:@19831.4]
  assign _T_25144 = _T_25143 | _T_25097; // @[Mux.scala 19:72:@19832.4]
  assign _T_25145 = _T_25144 | _T_25114; // @[Mux.scala 19:72:@19833.4]
  assign _T_25146 = _T_25145 | _T_25131; // @[Mux.scala 19:72:@19834.4]
  assign _T_25724 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0}; // @[Mux.scala 19:72:@20184.4]
  assign _T_25731 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8}; // @[Mux.scala 19:72:@20191.4]
  assign _T_25732 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,_T_25724}; // @[Mux.scala 19:72:@20192.4]
  assign _T_25734 = _T_2689 ? _T_25732 : 16'h0; // @[Mux.scala 19:72:@20193.4]
  assign _T_25741 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1}; // @[Mux.scala 19:72:@20200.4]
  assign _T_25748 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9}; // @[Mux.scala 19:72:@20207.4]
  assign _T_25749 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,_T_25741}; // @[Mux.scala 19:72:@20208.4]
  assign _T_25751 = _T_2690 ? _T_25749 : 16'h0; // @[Mux.scala 19:72:@20209.4]
  assign _T_25758 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2}; // @[Mux.scala 19:72:@20216.4]
  assign _T_25765 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10}; // @[Mux.scala 19:72:@20223.4]
  assign _T_25766 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,_T_25758}; // @[Mux.scala 19:72:@20224.4]
  assign _T_25768 = _T_2691 ? _T_25766 : 16'h0; // @[Mux.scala 19:72:@20225.4]
  assign _T_25775 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3}; // @[Mux.scala 19:72:@20232.4]
  assign _T_25782 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11}; // @[Mux.scala 19:72:@20239.4]
  assign _T_25783 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,_T_25775}; // @[Mux.scala 19:72:@20240.4]
  assign _T_25785 = _T_2692 ? _T_25783 : 16'h0; // @[Mux.scala 19:72:@20241.4]
  assign _T_25792 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4}; // @[Mux.scala 19:72:@20248.4]
  assign _T_25799 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12}; // @[Mux.scala 19:72:@20255.4]
  assign _T_25800 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,_T_25792}; // @[Mux.scala 19:72:@20256.4]
  assign _T_25802 = _T_2693 ? _T_25800 : 16'h0; // @[Mux.scala 19:72:@20257.4]
  assign _T_25809 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5}; // @[Mux.scala 19:72:@20264.4]
  assign _T_25816 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13}; // @[Mux.scala 19:72:@20271.4]
  assign _T_25817 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,_T_25809}; // @[Mux.scala 19:72:@20272.4]
  assign _T_25819 = _T_2694 ? _T_25817 : 16'h0; // @[Mux.scala 19:72:@20273.4]
  assign _T_25826 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6}; // @[Mux.scala 19:72:@20280.4]
  assign _T_25833 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14}; // @[Mux.scala 19:72:@20287.4]
  assign _T_25834 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,_T_25826}; // @[Mux.scala 19:72:@20288.4]
  assign _T_25836 = _T_2695 ? _T_25834 : 16'h0; // @[Mux.scala 19:72:@20289.4]
  assign _T_25843 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7}; // @[Mux.scala 19:72:@20296.4]
  assign _T_25850 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15}; // @[Mux.scala 19:72:@20303.4]
  assign _T_25851 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,_T_25843}; // @[Mux.scala 19:72:@20304.4]
  assign _T_25853 = _T_2696 ? _T_25851 : 16'h0; // @[Mux.scala 19:72:@20305.4]
  assign _T_25868 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,_T_25731}; // @[Mux.scala 19:72:@20320.4]
  assign _T_25870 = _T_2697 ? _T_25868 : 16'h0; // @[Mux.scala 19:72:@20321.4]
  assign _T_25885 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,_T_25748}; // @[Mux.scala 19:72:@20336.4]
  assign _T_25887 = _T_2698 ? _T_25885 : 16'h0; // @[Mux.scala 19:72:@20337.4]
  assign _T_25902 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,_T_25765}; // @[Mux.scala 19:72:@20352.4]
  assign _T_25904 = _T_2699 ? _T_25902 : 16'h0; // @[Mux.scala 19:72:@20353.4]
  assign _T_25919 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,_T_25782}; // @[Mux.scala 19:72:@20368.4]
  assign _T_25921 = _T_2700 ? _T_25919 : 16'h0; // @[Mux.scala 19:72:@20369.4]
  assign _T_25936 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,_T_25799}; // @[Mux.scala 19:72:@20384.4]
  assign _T_25938 = _T_2701 ? _T_25936 : 16'h0; // @[Mux.scala 19:72:@20385.4]
  assign _T_25953 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,_T_25816}; // @[Mux.scala 19:72:@20400.4]
  assign _T_25955 = _T_2702 ? _T_25953 : 16'h0; // @[Mux.scala 19:72:@20401.4]
  assign _T_25970 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,_T_25833}; // @[Mux.scala 19:72:@20416.4]
  assign _T_25972 = _T_2703 ? _T_25970 : 16'h0; // @[Mux.scala 19:72:@20417.4]
  assign _T_25987 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,_T_25850}; // @[Mux.scala 19:72:@20432.4]
  assign _T_25989 = _T_2704 ? _T_25987 : 16'h0; // @[Mux.scala 19:72:@20433.4]
  assign _T_25990 = _T_25734 | _T_25751; // @[Mux.scala 19:72:@20434.4]
  assign _T_25991 = _T_25990 | _T_25768; // @[Mux.scala 19:72:@20435.4]
  assign _T_25992 = _T_25991 | _T_25785; // @[Mux.scala 19:72:@20436.4]
  assign _T_25993 = _T_25992 | _T_25802; // @[Mux.scala 19:72:@20437.4]
  assign _T_25994 = _T_25993 | _T_25819; // @[Mux.scala 19:72:@20438.4]
  assign _T_25995 = _T_25994 | _T_25836; // @[Mux.scala 19:72:@20439.4]
  assign _T_25996 = _T_25995 | _T_25853; // @[Mux.scala 19:72:@20440.4]
  assign _T_25997 = _T_25996 | _T_25870; // @[Mux.scala 19:72:@20441.4]
  assign _T_25998 = _T_25997 | _T_25887; // @[Mux.scala 19:72:@20442.4]
  assign _T_25999 = _T_25998 | _T_25904; // @[Mux.scala 19:72:@20443.4]
  assign _T_26000 = _T_25999 | _T_25921; // @[Mux.scala 19:72:@20444.4]
  assign _T_26001 = _T_26000 | _T_25938; // @[Mux.scala 19:72:@20445.4]
  assign _T_26002 = _T_26001 | _T_25955; // @[Mux.scala 19:72:@20446.4]
  assign _T_26003 = _T_26002 | _T_25972; // @[Mux.scala 19:72:@20447.4]
  assign _T_26004 = _T_26003 | _T_25989; // @[Mux.scala 19:72:@20448.4]
  assign _T_26582 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0}; // @[Mux.scala 19:72:@20798.4]
  assign _T_26589 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8}; // @[Mux.scala 19:72:@20805.4]
  assign _T_26590 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,_T_26582}; // @[Mux.scala 19:72:@20806.4]
  assign _T_26592 = _T_2689 ? _T_26590 : 16'h0; // @[Mux.scala 19:72:@20807.4]
  assign _T_26599 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1}; // @[Mux.scala 19:72:@20814.4]
  assign _T_26606 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9}; // @[Mux.scala 19:72:@20821.4]
  assign _T_26607 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,_T_26599}; // @[Mux.scala 19:72:@20822.4]
  assign _T_26609 = _T_2690 ? _T_26607 : 16'h0; // @[Mux.scala 19:72:@20823.4]
  assign _T_26616 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2}; // @[Mux.scala 19:72:@20830.4]
  assign _T_26623 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10}; // @[Mux.scala 19:72:@20837.4]
  assign _T_26624 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,_T_26616}; // @[Mux.scala 19:72:@20838.4]
  assign _T_26626 = _T_2691 ? _T_26624 : 16'h0; // @[Mux.scala 19:72:@20839.4]
  assign _T_26633 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3}; // @[Mux.scala 19:72:@20846.4]
  assign _T_26640 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11}; // @[Mux.scala 19:72:@20853.4]
  assign _T_26641 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,_T_26633}; // @[Mux.scala 19:72:@20854.4]
  assign _T_26643 = _T_2692 ? _T_26641 : 16'h0; // @[Mux.scala 19:72:@20855.4]
  assign _T_26650 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4}; // @[Mux.scala 19:72:@20862.4]
  assign _T_26657 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12}; // @[Mux.scala 19:72:@20869.4]
  assign _T_26658 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,_T_26650}; // @[Mux.scala 19:72:@20870.4]
  assign _T_26660 = _T_2693 ? _T_26658 : 16'h0; // @[Mux.scala 19:72:@20871.4]
  assign _T_26667 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5}; // @[Mux.scala 19:72:@20878.4]
  assign _T_26674 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13}; // @[Mux.scala 19:72:@20885.4]
  assign _T_26675 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,_T_26667}; // @[Mux.scala 19:72:@20886.4]
  assign _T_26677 = _T_2694 ? _T_26675 : 16'h0; // @[Mux.scala 19:72:@20887.4]
  assign _T_26684 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6}; // @[Mux.scala 19:72:@20894.4]
  assign _T_26691 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14}; // @[Mux.scala 19:72:@20901.4]
  assign _T_26692 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,_T_26684}; // @[Mux.scala 19:72:@20902.4]
  assign _T_26694 = _T_2695 ? _T_26692 : 16'h0; // @[Mux.scala 19:72:@20903.4]
  assign _T_26701 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7}; // @[Mux.scala 19:72:@20910.4]
  assign _T_26708 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15}; // @[Mux.scala 19:72:@20917.4]
  assign _T_26709 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,_T_26701}; // @[Mux.scala 19:72:@20918.4]
  assign _T_26711 = _T_2696 ? _T_26709 : 16'h0; // @[Mux.scala 19:72:@20919.4]
  assign _T_26726 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,_T_26589}; // @[Mux.scala 19:72:@20934.4]
  assign _T_26728 = _T_2697 ? _T_26726 : 16'h0; // @[Mux.scala 19:72:@20935.4]
  assign _T_26743 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,_T_26606}; // @[Mux.scala 19:72:@20950.4]
  assign _T_26745 = _T_2698 ? _T_26743 : 16'h0; // @[Mux.scala 19:72:@20951.4]
  assign _T_26760 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,_T_26623}; // @[Mux.scala 19:72:@20966.4]
  assign _T_26762 = _T_2699 ? _T_26760 : 16'h0; // @[Mux.scala 19:72:@20967.4]
  assign _T_26777 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,_T_26640}; // @[Mux.scala 19:72:@20982.4]
  assign _T_26779 = _T_2700 ? _T_26777 : 16'h0; // @[Mux.scala 19:72:@20983.4]
  assign _T_26794 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,_T_26657}; // @[Mux.scala 19:72:@20998.4]
  assign _T_26796 = _T_2701 ? _T_26794 : 16'h0; // @[Mux.scala 19:72:@20999.4]
  assign _T_26811 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,_T_26674}; // @[Mux.scala 19:72:@21014.4]
  assign _T_26813 = _T_2702 ? _T_26811 : 16'h0; // @[Mux.scala 19:72:@21015.4]
  assign _T_26828 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,_T_26691}; // @[Mux.scala 19:72:@21030.4]
  assign _T_26830 = _T_2703 ? _T_26828 : 16'h0; // @[Mux.scala 19:72:@21031.4]
  assign _T_26845 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,_T_26708}; // @[Mux.scala 19:72:@21046.4]
  assign _T_26847 = _T_2704 ? _T_26845 : 16'h0; // @[Mux.scala 19:72:@21047.4]
  assign _T_26848 = _T_26592 | _T_26609; // @[Mux.scala 19:72:@21048.4]
  assign _T_26849 = _T_26848 | _T_26626; // @[Mux.scala 19:72:@21049.4]
  assign _T_26850 = _T_26849 | _T_26643; // @[Mux.scala 19:72:@21050.4]
  assign _T_26851 = _T_26850 | _T_26660; // @[Mux.scala 19:72:@21051.4]
  assign _T_26852 = _T_26851 | _T_26677; // @[Mux.scala 19:72:@21052.4]
  assign _T_26853 = _T_26852 | _T_26694; // @[Mux.scala 19:72:@21053.4]
  assign _T_26854 = _T_26853 | _T_26711; // @[Mux.scala 19:72:@21054.4]
  assign _T_26855 = _T_26854 | _T_26728; // @[Mux.scala 19:72:@21055.4]
  assign _T_26856 = _T_26855 | _T_26745; // @[Mux.scala 19:72:@21056.4]
  assign _T_26857 = _T_26856 | _T_26762; // @[Mux.scala 19:72:@21057.4]
  assign _T_26858 = _T_26857 | _T_26779; // @[Mux.scala 19:72:@21058.4]
  assign _T_26859 = _T_26858 | _T_26796; // @[Mux.scala 19:72:@21059.4]
  assign _T_26860 = _T_26859 | _T_26813; // @[Mux.scala 19:72:@21060.4]
  assign _T_26861 = _T_26860 | _T_26830; // @[Mux.scala 19:72:@21061.4]
  assign _T_26862 = _T_26861 | _T_26847; // @[Mux.scala 19:72:@21062.4]
  assign _T_27440 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0}; // @[Mux.scala 19:72:@21412.4]
  assign _T_27447 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8}; // @[Mux.scala 19:72:@21419.4]
  assign _T_27448 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,_T_27440}; // @[Mux.scala 19:72:@21420.4]
  assign _T_27450 = _T_2689 ? _T_27448 : 16'h0; // @[Mux.scala 19:72:@21421.4]
  assign _T_27457 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1}; // @[Mux.scala 19:72:@21428.4]
  assign _T_27464 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9}; // @[Mux.scala 19:72:@21435.4]
  assign _T_27465 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,_T_27457}; // @[Mux.scala 19:72:@21436.4]
  assign _T_27467 = _T_2690 ? _T_27465 : 16'h0; // @[Mux.scala 19:72:@21437.4]
  assign _T_27474 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2}; // @[Mux.scala 19:72:@21444.4]
  assign _T_27481 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10}; // @[Mux.scala 19:72:@21451.4]
  assign _T_27482 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,_T_27474}; // @[Mux.scala 19:72:@21452.4]
  assign _T_27484 = _T_2691 ? _T_27482 : 16'h0; // @[Mux.scala 19:72:@21453.4]
  assign _T_27491 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3}; // @[Mux.scala 19:72:@21460.4]
  assign _T_27498 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11}; // @[Mux.scala 19:72:@21467.4]
  assign _T_27499 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,_T_27491}; // @[Mux.scala 19:72:@21468.4]
  assign _T_27501 = _T_2692 ? _T_27499 : 16'h0; // @[Mux.scala 19:72:@21469.4]
  assign _T_27508 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4}; // @[Mux.scala 19:72:@21476.4]
  assign _T_27515 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12}; // @[Mux.scala 19:72:@21483.4]
  assign _T_27516 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,_T_27508}; // @[Mux.scala 19:72:@21484.4]
  assign _T_27518 = _T_2693 ? _T_27516 : 16'h0; // @[Mux.scala 19:72:@21485.4]
  assign _T_27525 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5}; // @[Mux.scala 19:72:@21492.4]
  assign _T_27532 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13}; // @[Mux.scala 19:72:@21499.4]
  assign _T_27533 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,_T_27525}; // @[Mux.scala 19:72:@21500.4]
  assign _T_27535 = _T_2694 ? _T_27533 : 16'h0; // @[Mux.scala 19:72:@21501.4]
  assign _T_27542 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6}; // @[Mux.scala 19:72:@21508.4]
  assign _T_27549 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14}; // @[Mux.scala 19:72:@21515.4]
  assign _T_27550 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,_T_27542}; // @[Mux.scala 19:72:@21516.4]
  assign _T_27552 = _T_2695 ? _T_27550 : 16'h0; // @[Mux.scala 19:72:@21517.4]
  assign _T_27559 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7}; // @[Mux.scala 19:72:@21524.4]
  assign _T_27566 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15}; // @[Mux.scala 19:72:@21531.4]
  assign _T_27567 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,_T_27559}; // @[Mux.scala 19:72:@21532.4]
  assign _T_27569 = _T_2696 ? _T_27567 : 16'h0; // @[Mux.scala 19:72:@21533.4]
  assign _T_27584 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,_T_27447}; // @[Mux.scala 19:72:@21548.4]
  assign _T_27586 = _T_2697 ? _T_27584 : 16'h0; // @[Mux.scala 19:72:@21549.4]
  assign _T_27601 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,_T_27464}; // @[Mux.scala 19:72:@21564.4]
  assign _T_27603 = _T_2698 ? _T_27601 : 16'h0; // @[Mux.scala 19:72:@21565.4]
  assign _T_27618 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,_T_27481}; // @[Mux.scala 19:72:@21580.4]
  assign _T_27620 = _T_2699 ? _T_27618 : 16'h0; // @[Mux.scala 19:72:@21581.4]
  assign _T_27635 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,_T_27498}; // @[Mux.scala 19:72:@21596.4]
  assign _T_27637 = _T_2700 ? _T_27635 : 16'h0; // @[Mux.scala 19:72:@21597.4]
  assign _T_27652 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,_T_27515}; // @[Mux.scala 19:72:@21612.4]
  assign _T_27654 = _T_2701 ? _T_27652 : 16'h0; // @[Mux.scala 19:72:@21613.4]
  assign _T_27669 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,_T_27532}; // @[Mux.scala 19:72:@21628.4]
  assign _T_27671 = _T_2702 ? _T_27669 : 16'h0; // @[Mux.scala 19:72:@21629.4]
  assign _T_27686 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,_T_27549}; // @[Mux.scala 19:72:@21644.4]
  assign _T_27688 = _T_2703 ? _T_27686 : 16'h0; // @[Mux.scala 19:72:@21645.4]
  assign _T_27703 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,_T_27566}; // @[Mux.scala 19:72:@21660.4]
  assign _T_27705 = _T_2704 ? _T_27703 : 16'h0; // @[Mux.scala 19:72:@21661.4]
  assign _T_27706 = _T_27450 | _T_27467; // @[Mux.scala 19:72:@21662.4]
  assign _T_27707 = _T_27706 | _T_27484; // @[Mux.scala 19:72:@21663.4]
  assign _T_27708 = _T_27707 | _T_27501; // @[Mux.scala 19:72:@21664.4]
  assign _T_27709 = _T_27708 | _T_27518; // @[Mux.scala 19:72:@21665.4]
  assign _T_27710 = _T_27709 | _T_27535; // @[Mux.scala 19:72:@21666.4]
  assign _T_27711 = _T_27710 | _T_27552; // @[Mux.scala 19:72:@21667.4]
  assign _T_27712 = _T_27711 | _T_27569; // @[Mux.scala 19:72:@21668.4]
  assign _T_27713 = _T_27712 | _T_27586; // @[Mux.scala 19:72:@21669.4]
  assign _T_27714 = _T_27713 | _T_27603; // @[Mux.scala 19:72:@21670.4]
  assign _T_27715 = _T_27714 | _T_27620; // @[Mux.scala 19:72:@21671.4]
  assign _T_27716 = _T_27715 | _T_27637; // @[Mux.scala 19:72:@21672.4]
  assign _T_27717 = _T_27716 | _T_27654; // @[Mux.scala 19:72:@21673.4]
  assign _T_27718 = _T_27717 | _T_27671; // @[Mux.scala 19:72:@21674.4]
  assign _T_27719 = _T_27718 | _T_27688; // @[Mux.scala 19:72:@21675.4]
  assign _T_27720 = _T_27719 | _T_27705; // @[Mux.scala 19:72:@21676.4]
  assign _T_28298 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0}; // @[Mux.scala 19:72:@22026.4]
  assign _T_28305 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8}; // @[Mux.scala 19:72:@22033.4]
  assign _T_28306 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,_T_28298}; // @[Mux.scala 19:72:@22034.4]
  assign _T_28308 = _T_2689 ? _T_28306 : 16'h0; // @[Mux.scala 19:72:@22035.4]
  assign _T_28315 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1}; // @[Mux.scala 19:72:@22042.4]
  assign _T_28322 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9}; // @[Mux.scala 19:72:@22049.4]
  assign _T_28323 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,_T_28315}; // @[Mux.scala 19:72:@22050.4]
  assign _T_28325 = _T_2690 ? _T_28323 : 16'h0; // @[Mux.scala 19:72:@22051.4]
  assign _T_28332 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2}; // @[Mux.scala 19:72:@22058.4]
  assign _T_28339 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10}; // @[Mux.scala 19:72:@22065.4]
  assign _T_28340 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,_T_28332}; // @[Mux.scala 19:72:@22066.4]
  assign _T_28342 = _T_2691 ? _T_28340 : 16'h0; // @[Mux.scala 19:72:@22067.4]
  assign _T_28349 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3}; // @[Mux.scala 19:72:@22074.4]
  assign _T_28356 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11}; // @[Mux.scala 19:72:@22081.4]
  assign _T_28357 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,_T_28349}; // @[Mux.scala 19:72:@22082.4]
  assign _T_28359 = _T_2692 ? _T_28357 : 16'h0; // @[Mux.scala 19:72:@22083.4]
  assign _T_28366 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4}; // @[Mux.scala 19:72:@22090.4]
  assign _T_28373 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12}; // @[Mux.scala 19:72:@22097.4]
  assign _T_28374 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,_T_28366}; // @[Mux.scala 19:72:@22098.4]
  assign _T_28376 = _T_2693 ? _T_28374 : 16'h0; // @[Mux.scala 19:72:@22099.4]
  assign _T_28383 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5}; // @[Mux.scala 19:72:@22106.4]
  assign _T_28390 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13}; // @[Mux.scala 19:72:@22113.4]
  assign _T_28391 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,_T_28383}; // @[Mux.scala 19:72:@22114.4]
  assign _T_28393 = _T_2694 ? _T_28391 : 16'h0; // @[Mux.scala 19:72:@22115.4]
  assign _T_28400 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6}; // @[Mux.scala 19:72:@22122.4]
  assign _T_28407 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14}; // @[Mux.scala 19:72:@22129.4]
  assign _T_28408 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,_T_28400}; // @[Mux.scala 19:72:@22130.4]
  assign _T_28410 = _T_2695 ? _T_28408 : 16'h0; // @[Mux.scala 19:72:@22131.4]
  assign _T_28417 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7}; // @[Mux.scala 19:72:@22138.4]
  assign _T_28424 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15}; // @[Mux.scala 19:72:@22145.4]
  assign _T_28425 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,_T_28417}; // @[Mux.scala 19:72:@22146.4]
  assign _T_28427 = _T_2696 ? _T_28425 : 16'h0; // @[Mux.scala 19:72:@22147.4]
  assign _T_28442 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,_T_28305}; // @[Mux.scala 19:72:@22162.4]
  assign _T_28444 = _T_2697 ? _T_28442 : 16'h0; // @[Mux.scala 19:72:@22163.4]
  assign _T_28459 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,_T_28322}; // @[Mux.scala 19:72:@22178.4]
  assign _T_28461 = _T_2698 ? _T_28459 : 16'h0; // @[Mux.scala 19:72:@22179.4]
  assign _T_28476 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,_T_28339}; // @[Mux.scala 19:72:@22194.4]
  assign _T_28478 = _T_2699 ? _T_28476 : 16'h0; // @[Mux.scala 19:72:@22195.4]
  assign _T_28493 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,_T_28356}; // @[Mux.scala 19:72:@22210.4]
  assign _T_28495 = _T_2700 ? _T_28493 : 16'h0; // @[Mux.scala 19:72:@22211.4]
  assign _T_28510 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,_T_28373}; // @[Mux.scala 19:72:@22226.4]
  assign _T_28512 = _T_2701 ? _T_28510 : 16'h0; // @[Mux.scala 19:72:@22227.4]
  assign _T_28527 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,_T_28390}; // @[Mux.scala 19:72:@22242.4]
  assign _T_28529 = _T_2702 ? _T_28527 : 16'h0; // @[Mux.scala 19:72:@22243.4]
  assign _T_28544 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,_T_28407}; // @[Mux.scala 19:72:@22258.4]
  assign _T_28546 = _T_2703 ? _T_28544 : 16'h0; // @[Mux.scala 19:72:@22259.4]
  assign _T_28561 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,_T_28424}; // @[Mux.scala 19:72:@22274.4]
  assign _T_28563 = _T_2704 ? _T_28561 : 16'h0; // @[Mux.scala 19:72:@22275.4]
  assign _T_28564 = _T_28308 | _T_28325; // @[Mux.scala 19:72:@22276.4]
  assign _T_28565 = _T_28564 | _T_28342; // @[Mux.scala 19:72:@22277.4]
  assign _T_28566 = _T_28565 | _T_28359; // @[Mux.scala 19:72:@22278.4]
  assign _T_28567 = _T_28566 | _T_28376; // @[Mux.scala 19:72:@22279.4]
  assign _T_28568 = _T_28567 | _T_28393; // @[Mux.scala 19:72:@22280.4]
  assign _T_28569 = _T_28568 | _T_28410; // @[Mux.scala 19:72:@22281.4]
  assign _T_28570 = _T_28569 | _T_28427; // @[Mux.scala 19:72:@22282.4]
  assign _T_28571 = _T_28570 | _T_28444; // @[Mux.scala 19:72:@22283.4]
  assign _T_28572 = _T_28571 | _T_28461; // @[Mux.scala 19:72:@22284.4]
  assign _T_28573 = _T_28572 | _T_28478; // @[Mux.scala 19:72:@22285.4]
  assign _T_28574 = _T_28573 | _T_28495; // @[Mux.scala 19:72:@22286.4]
  assign _T_28575 = _T_28574 | _T_28512; // @[Mux.scala 19:72:@22287.4]
  assign _T_28576 = _T_28575 | _T_28529; // @[Mux.scala 19:72:@22288.4]
  assign _T_28577 = _T_28576 | _T_28546; // @[Mux.scala 19:72:@22289.4]
  assign _T_28578 = _T_28577 | _T_28563; // @[Mux.scala 19:72:@22290.4]
  assign _T_29156 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0}; // @[Mux.scala 19:72:@22640.4]
  assign _T_29163 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8}; // @[Mux.scala 19:72:@22647.4]
  assign _T_29164 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,_T_29156}; // @[Mux.scala 19:72:@22648.4]
  assign _T_29166 = _T_2689 ? _T_29164 : 16'h0; // @[Mux.scala 19:72:@22649.4]
  assign _T_29173 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1}; // @[Mux.scala 19:72:@22656.4]
  assign _T_29180 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9}; // @[Mux.scala 19:72:@22663.4]
  assign _T_29181 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,_T_29173}; // @[Mux.scala 19:72:@22664.4]
  assign _T_29183 = _T_2690 ? _T_29181 : 16'h0; // @[Mux.scala 19:72:@22665.4]
  assign _T_29190 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2}; // @[Mux.scala 19:72:@22672.4]
  assign _T_29197 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10}; // @[Mux.scala 19:72:@22679.4]
  assign _T_29198 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,_T_29190}; // @[Mux.scala 19:72:@22680.4]
  assign _T_29200 = _T_2691 ? _T_29198 : 16'h0; // @[Mux.scala 19:72:@22681.4]
  assign _T_29207 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3}; // @[Mux.scala 19:72:@22688.4]
  assign _T_29214 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11}; // @[Mux.scala 19:72:@22695.4]
  assign _T_29215 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,_T_29207}; // @[Mux.scala 19:72:@22696.4]
  assign _T_29217 = _T_2692 ? _T_29215 : 16'h0; // @[Mux.scala 19:72:@22697.4]
  assign _T_29224 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4}; // @[Mux.scala 19:72:@22704.4]
  assign _T_29231 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12}; // @[Mux.scala 19:72:@22711.4]
  assign _T_29232 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,_T_29224}; // @[Mux.scala 19:72:@22712.4]
  assign _T_29234 = _T_2693 ? _T_29232 : 16'h0; // @[Mux.scala 19:72:@22713.4]
  assign _T_29241 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5}; // @[Mux.scala 19:72:@22720.4]
  assign _T_29248 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13}; // @[Mux.scala 19:72:@22727.4]
  assign _T_29249 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,_T_29241}; // @[Mux.scala 19:72:@22728.4]
  assign _T_29251 = _T_2694 ? _T_29249 : 16'h0; // @[Mux.scala 19:72:@22729.4]
  assign _T_29258 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6}; // @[Mux.scala 19:72:@22736.4]
  assign _T_29265 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14}; // @[Mux.scala 19:72:@22743.4]
  assign _T_29266 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,_T_29258}; // @[Mux.scala 19:72:@22744.4]
  assign _T_29268 = _T_2695 ? _T_29266 : 16'h0; // @[Mux.scala 19:72:@22745.4]
  assign _T_29275 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7}; // @[Mux.scala 19:72:@22752.4]
  assign _T_29282 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15}; // @[Mux.scala 19:72:@22759.4]
  assign _T_29283 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,_T_29275}; // @[Mux.scala 19:72:@22760.4]
  assign _T_29285 = _T_2696 ? _T_29283 : 16'h0; // @[Mux.scala 19:72:@22761.4]
  assign _T_29300 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,_T_29163}; // @[Mux.scala 19:72:@22776.4]
  assign _T_29302 = _T_2697 ? _T_29300 : 16'h0; // @[Mux.scala 19:72:@22777.4]
  assign _T_29317 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,_T_29180}; // @[Mux.scala 19:72:@22792.4]
  assign _T_29319 = _T_2698 ? _T_29317 : 16'h0; // @[Mux.scala 19:72:@22793.4]
  assign _T_29334 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,_T_29197}; // @[Mux.scala 19:72:@22808.4]
  assign _T_29336 = _T_2699 ? _T_29334 : 16'h0; // @[Mux.scala 19:72:@22809.4]
  assign _T_29351 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,_T_29214}; // @[Mux.scala 19:72:@22824.4]
  assign _T_29353 = _T_2700 ? _T_29351 : 16'h0; // @[Mux.scala 19:72:@22825.4]
  assign _T_29368 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,_T_29231}; // @[Mux.scala 19:72:@22840.4]
  assign _T_29370 = _T_2701 ? _T_29368 : 16'h0; // @[Mux.scala 19:72:@22841.4]
  assign _T_29385 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,_T_29248}; // @[Mux.scala 19:72:@22856.4]
  assign _T_29387 = _T_2702 ? _T_29385 : 16'h0; // @[Mux.scala 19:72:@22857.4]
  assign _T_29402 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,_T_29265}; // @[Mux.scala 19:72:@22872.4]
  assign _T_29404 = _T_2703 ? _T_29402 : 16'h0; // @[Mux.scala 19:72:@22873.4]
  assign _T_29419 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,_T_29282}; // @[Mux.scala 19:72:@22888.4]
  assign _T_29421 = _T_2704 ? _T_29419 : 16'h0; // @[Mux.scala 19:72:@22889.4]
  assign _T_29422 = _T_29166 | _T_29183; // @[Mux.scala 19:72:@22890.4]
  assign _T_29423 = _T_29422 | _T_29200; // @[Mux.scala 19:72:@22891.4]
  assign _T_29424 = _T_29423 | _T_29217; // @[Mux.scala 19:72:@22892.4]
  assign _T_29425 = _T_29424 | _T_29234; // @[Mux.scala 19:72:@22893.4]
  assign _T_29426 = _T_29425 | _T_29251; // @[Mux.scala 19:72:@22894.4]
  assign _T_29427 = _T_29426 | _T_29268; // @[Mux.scala 19:72:@22895.4]
  assign _T_29428 = _T_29427 | _T_29285; // @[Mux.scala 19:72:@22896.4]
  assign _T_29429 = _T_29428 | _T_29302; // @[Mux.scala 19:72:@22897.4]
  assign _T_29430 = _T_29429 | _T_29319; // @[Mux.scala 19:72:@22898.4]
  assign _T_29431 = _T_29430 | _T_29336; // @[Mux.scala 19:72:@22899.4]
  assign _T_29432 = _T_29431 | _T_29353; // @[Mux.scala 19:72:@22900.4]
  assign _T_29433 = _T_29432 | _T_29370; // @[Mux.scala 19:72:@22901.4]
  assign _T_29434 = _T_29433 | _T_29387; // @[Mux.scala 19:72:@22902.4]
  assign _T_29435 = _T_29434 | _T_29404; // @[Mux.scala 19:72:@22903.4]
  assign _T_29436 = _T_29435 | _T_29421; // @[Mux.scala 19:72:@22904.4]
  assign _T_30014 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0}; // @[Mux.scala 19:72:@23254.4]
  assign _T_30021 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8}; // @[Mux.scala 19:72:@23261.4]
  assign _T_30022 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,_T_30014}; // @[Mux.scala 19:72:@23262.4]
  assign _T_30024 = _T_2689 ? _T_30022 : 16'h0; // @[Mux.scala 19:72:@23263.4]
  assign _T_30031 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1}; // @[Mux.scala 19:72:@23270.4]
  assign _T_30038 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9}; // @[Mux.scala 19:72:@23277.4]
  assign _T_30039 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,_T_30031}; // @[Mux.scala 19:72:@23278.4]
  assign _T_30041 = _T_2690 ? _T_30039 : 16'h0; // @[Mux.scala 19:72:@23279.4]
  assign _T_30048 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2}; // @[Mux.scala 19:72:@23286.4]
  assign _T_30055 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10}; // @[Mux.scala 19:72:@23293.4]
  assign _T_30056 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,_T_30048}; // @[Mux.scala 19:72:@23294.4]
  assign _T_30058 = _T_2691 ? _T_30056 : 16'h0; // @[Mux.scala 19:72:@23295.4]
  assign _T_30065 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3}; // @[Mux.scala 19:72:@23302.4]
  assign _T_30072 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11}; // @[Mux.scala 19:72:@23309.4]
  assign _T_30073 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,_T_30065}; // @[Mux.scala 19:72:@23310.4]
  assign _T_30075 = _T_2692 ? _T_30073 : 16'h0; // @[Mux.scala 19:72:@23311.4]
  assign _T_30082 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4}; // @[Mux.scala 19:72:@23318.4]
  assign _T_30089 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12}; // @[Mux.scala 19:72:@23325.4]
  assign _T_30090 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,_T_30082}; // @[Mux.scala 19:72:@23326.4]
  assign _T_30092 = _T_2693 ? _T_30090 : 16'h0; // @[Mux.scala 19:72:@23327.4]
  assign _T_30099 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5}; // @[Mux.scala 19:72:@23334.4]
  assign _T_30106 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13}; // @[Mux.scala 19:72:@23341.4]
  assign _T_30107 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,_T_30099}; // @[Mux.scala 19:72:@23342.4]
  assign _T_30109 = _T_2694 ? _T_30107 : 16'h0; // @[Mux.scala 19:72:@23343.4]
  assign _T_30116 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6}; // @[Mux.scala 19:72:@23350.4]
  assign _T_30123 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14}; // @[Mux.scala 19:72:@23357.4]
  assign _T_30124 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,_T_30116}; // @[Mux.scala 19:72:@23358.4]
  assign _T_30126 = _T_2695 ? _T_30124 : 16'h0; // @[Mux.scala 19:72:@23359.4]
  assign _T_30133 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7}; // @[Mux.scala 19:72:@23366.4]
  assign _T_30140 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15}; // @[Mux.scala 19:72:@23373.4]
  assign _T_30141 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,_T_30133}; // @[Mux.scala 19:72:@23374.4]
  assign _T_30143 = _T_2696 ? _T_30141 : 16'h0; // @[Mux.scala 19:72:@23375.4]
  assign _T_30158 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,_T_30021}; // @[Mux.scala 19:72:@23390.4]
  assign _T_30160 = _T_2697 ? _T_30158 : 16'h0; // @[Mux.scala 19:72:@23391.4]
  assign _T_30175 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,_T_30038}; // @[Mux.scala 19:72:@23406.4]
  assign _T_30177 = _T_2698 ? _T_30175 : 16'h0; // @[Mux.scala 19:72:@23407.4]
  assign _T_30192 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,_T_30055}; // @[Mux.scala 19:72:@23422.4]
  assign _T_30194 = _T_2699 ? _T_30192 : 16'h0; // @[Mux.scala 19:72:@23423.4]
  assign _T_30209 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,_T_30072}; // @[Mux.scala 19:72:@23438.4]
  assign _T_30211 = _T_2700 ? _T_30209 : 16'h0; // @[Mux.scala 19:72:@23439.4]
  assign _T_30226 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,_T_30089}; // @[Mux.scala 19:72:@23454.4]
  assign _T_30228 = _T_2701 ? _T_30226 : 16'h0; // @[Mux.scala 19:72:@23455.4]
  assign _T_30243 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,_T_30106}; // @[Mux.scala 19:72:@23470.4]
  assign _T_30245 = _T_2702 ? _T_30243 : 16'h0; // @[Mux.scala 19:72:@23471.4]
  assign _T_30260 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,_T_30123}; // @[Mux.scala 19:72:@23486.4]
  assign _T_30262 = _T_2703 ? _T_30260 : 16'h0; // @[Mux.scala 19:72:@23487.4]
  assign _T_30277 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,_T_30140}; // @[Mux.scala 19:72:@23502.4]
  assign _T_30279 = _T_2704 ? _T_30277 : 16'h0; // @[Mux.scala 19:72:@23503.4]
  assign _T_30280 = _T_30024 | _T_30041; // @[Mux.scala 19:72:@23504.4]
  assign _T_30281 = _T_30280 | _T_30058; // @[Mux.scala 19:72:@23505.4]
  assign _T_30282 = _T_30281 | _T_30075; // @[Mux.scala 19:72:@23506.4]
  assign _T_30283 = _T_30282 | _T_30092; // @[Mux.scala 19:72:@23507.4]
  assign _T_30284 = _T_30283 | _T_30109; // @[Mux.scala 19:72:@23508.4]
  assign _T_30285 = _T_30284 | _T_30126; // @[Mux.scala 19:72:@23509.4]
  assign _T_30286 = _T_30285 | _T_30143; // @[Mux.scala 19:72:@23510.4]
  assign _T_30287 = _T_30286 | _T_30160; // @[Mux.scala 19:72:@23511.4]
  assign _T_30288 = _T_30287 | _T_30177; // @[Mux.scala 19:72:@23512.4]
  assign _T_30289 = _T_30288 | _T_30194; // @[Mux.scala 19:72:@23513.4]
  assign _T_30290 = _T_30289 | _T_30211; // @[Mux.scala 19:72:@23514.4]
  assign _T_30291 = _T_30290 | _T_30228; // @[Mux.scala 19:72:@23515.4]
  assign _T_30292 = _T_30291 | _T_30245; // @[Mux.scala 19:72:@23516.4]
  assign _T_30293 = _T_30292 | _T_30262; // @[Mux.scala 19:72:@23517.4]
  assign _T_30294 = _T_30293 | _T_30279; // @[Mux.scala 19:72:@23518.4]
  assign _T_30872 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0}; // @[Mux.scala 19:72:@23868.4]
  assign _T_30879 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8}; // @[Mux.scala 19:72:@23875.4]
  assign _T_30880 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,_T_30872}; // @[Mux.scala 19:72:@23876.4]
  assign _T_30882 = _T_2689 ? _T_30880 : 16'h0; // @[Mux.scala 19:72:@23877.4]
  assign _T_30889 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1}; // @[Mux.scala 19:72:@23884.4]
  assign _T_30896 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9}; // @[Mux.scala 19:72:@23891.4]
  assign _T_30897 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,_T_30889}; // @[Mux.scala 19:72:@23892.4]
  assign _T_30899 = _T_2690 ? _T_30897 : 16'h0; // @[Mux.scala 19:72:@23893.4]
  assign _T_30906 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2}; // @[Mux.scala 19:72:@23900.4]
  assign _T_30913 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10}; // @[Mux.scala 19:72:@23907.4]
  assign _T_30914 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,_T_30906}; // @[Mux.scala 19:72:@23908.4]
  assign _T_30916 = _T_2691 ? _T_30914 : 16'h0; // @[Mux.scala 19:72:@23909.4]
  assign _T_30923 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3}; // @[Mux.scala 19:72:@23916.4]
  assign _T_30930 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11}; // @[Mux.scala 19:72:@23923.4]
  assign _T_30931 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,_T_30923}; // @[Mux.scala 19:72:@23924.4]
  assign _T_30933 = _T_2692 ? _T_30931 : 16'h0; // @[Mux.scala 19:72:@23925.4]
  assign _T_30940 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4}; // @[Mux.scala 19:72:@23932.4]
  assign _T_30947 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12}; // @[Mux.scala 19:72:@23939.4]
  assign _T_30948 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,_T_30940}; // @[Mux.scala 19:72:@23940.4]
  assign _T_30950 = _T_2693 ? _T_30948 : 16'h0; // @[Mux.scala 19:72:@23941.4]
  assign _T_30957 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5}; // @[Mux.scala 19:72:@23948.4]
  assign _T_30964 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13}; // @[Mux.scala 19:72:@23955.4]
  assign _T_30965 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,_T_30957}; // @[Mux.scala 19:72:@23956.4]
  assign _T_30967 = _T_2694 ? _T_30965 : 16'h0; // @[Mux.scala 19:72:@23957.4]
  assign _T_30974 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6}; // @[Mux.scala 19:72:@23964.4]
  assign _T_30981 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14}; // @[Mux.scala 19:72:@23971.4]
  assign _T_30982 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,_T_30974}; // @[Mux.scala 19:72:@23972.4]
  assign _T_30984 = _T_2695 ? _T_30982 : 16'h0; // @[Mux.scala 19:72:@23973.4]
  assign _T_30991 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7}; // @[Mux.scala 19:72:@23980.4]
  assign _T_30998 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15}; // @[Mux.scala 19:72:@23987.4]
  assign _T_30999 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,_T_30991}; // @[Mux.scala 19:72:@23988.4]
  assign _T_31001 = _T_2696 ? _T_30999 : 16'h0; // @[Mux.scala 19:72:@23989.4]
  assign _T_31016 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,_T_30879}; // @[Mux.scala 19:72:@24004.4]
  assign _T_31018 = _T_2697 ? _T_31016 : 16'h0; // @[Mux.scala 19:72:@24005.4]
  assign _T_31033 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,_T_30896}; // @[Mux.scala 19:72:@24020.4]
  assign _T_31035 = _T_2698 ? _T_31033 : 16'h0; // @[Mux.scala 19:72:@24021.4]
  assign _T_31050 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,_T_30913}; // @[Mux.scala 19:72:@24036.4]
  assign _T_31052 = _T_2699 ? _T_31050 : 16'h0; // @[Mux.scala 19:72:@24037.4]
  assign _T_31067 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,_T_30930}; // @[Mux.scala 19:72:@24052.4]
  assign _T_31069 = _T_2700 ? _T_31067 : 16'h0; // @[Mux.scala 19:72:@24053.4]
  assign _T_31084 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,_T_30947}; // @[Mux.scala 19:72:@24068.4]
  assign _T_31086 = _T_2701 ? _T_31084 : 16'h0; // @[Mux.scala 19:72:@24069.4]
  assign _T_31101 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,_T_30964}; // @[Mux.scala 19:72:@24084.4]
  assign _T_31103 = _T_2702 ? _T_31101 : 16'h0; // @[Mux.scala 19:72:@24085.4]
  assign _T_31118 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,_T_30981}; // @[Mux.scala 19:72:@24100.4]
  assign _T_31120 = _T_2703 ? _T_31118 : 16'h0; // @[Mux.scala 19:72:@24101.4]
  assign _T_31135 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,_T_30998}; // @[Mux.scala 19:72:@24116.4]
  assign _T_31137 = _T_2704 ? _T_31135 : 16'h0; // @[Mux.scala 19:72:@24117.4]
  assign _T_31138 = _T_30882 | _T_30899; // @[Mux.scala 19:72:@24118.4]
  assign _T_31139 = _T_31138 | _T_30916; // @[Mux.scala 19:72:@24119.4]
  assign _T_31140 = _T_31139 | _T_30933; // @[Mux.scala 19:72:@24120.4]
  assign _T_31141 = _T_31140 | _T_30950; // @[Mux.scala 19:72:@24121.4]
  assign _T_31142 = _T_31141 | _T_30967; // @[Mux.scala 19:72:@24122.4]
  assign _T_31143 = _T_31142 | _T_30984; // @[Mux.scala 19:72:@24123.4]
  assign _T_31144 = _T_31143 | _T_31001; // @[Mux.scala 19:72:@24124.4]
  assign _T_31145 = _T_31144 | _T_31018; // @[Mux.scala 19:72:@24125.4]
  assign _T_31146 = _T_31145 | _T_31035; // @[Mux.scala 19:72:@24126.4]
  assign _T_31147 = _T_31146 | _T_31052; // @[Mux.scala 19:72:@24127.4]
  assign _T_31148 = _T_31147 | _T_31069; // @[Mux.scala 19:72:@24128.4]
  assign _T_31149 = _T_31148 | _T_31086; // @[Mux.scala 19:72:@24129.4]
  assign _T_31150 = _T_31149 | _T_31103; // @[Mux.scala 19:72:@24130.4]
  assign _T_31151 = _T_31150 | _T_31120; // @[Mux.scala 19:72:@24131.4]
  assign _T_31152 = _T_31151 | _T_31137; // @[Mux.scala 19:72:@24132.4]
  assign _T_52326 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@24996.4]
  assign _T_52333 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8}; // @[Mux.scala 19:72:@25003.4]
  assign _T_52334 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,_T_52326}; // @[Mux.scala 19:72:@25004.4]
  assign _T_52336 = _T_2689 ? _T_52334 : 16'h0; // @[Mux.scala 19:72:@25005.4]
  assign _T_52343 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@25012.4]
  assign _T_52350 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9}; // @[Mux.scala 19:72:@25019.4]
  assign _T_52351 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,_T_52343}; // @[Mux.scala 19:72:@25020.4]
  assign _T_52353 = _T_2690 ? _T_52351 : 16'h0; // @[Mux.scala 19:72:@25021.4]
  assign _T_52360 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@25028.4]
  assign _T_52367 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10}; // @[Mux.scala 19:72:@25035.4]
  assign _T_52368 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,_T_52360}; // @[Mux.scala 19:72:@25036.4]
  assign _T_52370 = _T_2691 ? _T_52368 : 16'h0; // @[Mux.scala 19:72:@25037.4]
  assign _T_52377 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@25044.4]
  assign _T_52384 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11}; // @[Mux.scala 19:72:@25051.4]
  assign _T_52385 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,_T_52377}; // @[Mux.scala 19:72:@25052.4]
  assign _T_52387 = _T_2692 ? _T_52385 : 16'h0; // @[Mux.scala 19:72:@25053.4]
  assign _T_52394 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@25060.4]
  assign _T_52401 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12}; // @[Mux.scala 19:72:@25067.4]
  assign _T_52402 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,_T_52394}; // @[Mux.scala 19:72:@25068.4]
  assign _T_52404 = _T_2693 ? _T_52402 : 16'h0; // @[Mux.scala 19:72:@25069.4]
  assign _T_52411 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@25076.4]
  assign _T_52418 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13}; // @[Mux.scala 19:72:@25083.4]
  assign _T_52419 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,_T_52411}; // @[Mux.scala 19:72:@25084.4]
  assign _T_52421 = _T_2694 ? _T_52419 : 16'h0; // @[Mux.scala 19:72:@25085.4]
  assign _T_52428 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@25092.4]
  assign _T_52435 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14}; // @[Mux.scala 19:72:@25099.4]
  assign _T_52436 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,_T_52428}; // @[Mux.scala 19:72:@25100.4]
  assign _T_52438 = _T_2695 ? _T_52436 : 16'h0; // @[Mux.scala 19:72:@25101.4]
  assign _T_52445 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@25108.4]
  assign _T_52452 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15}; // @[Mux.scala 19:72:@25115.4]
  assign _T_52453 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,_T_52445}; // @[Mux.scala 19:72:@25116.4]
  assign _T_52455 = _T_2696 ? _T_52453 : 16'h0; // @[Mux.scala 19:72:@25117.4]
  assign _T_52470 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,_T_52333}; // @[Mux.scala 19:72:@25132.4]
  assign _T_52472 = _T_2697 ? _T_52470 : 16'h0; // @[Mux.scala 19:72:@25133.4]
  assign _T_52487 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,_T_52350}; // @[Mux.scala 19:72:@25148.4]
  assign _T_52489 = _T_2698 ? _T_52487 : 16'h0; // @[Mux.scala 19:72:@25149.4]
  assign _T_52504 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,_T_52367}; // @[Mux.scala 19:72:@25164.4]
  assign _T_52506 = _T_2699 ? _T_52504 : 16'h0; // @[Mux.scala 19:72:@25165.4]
  assign _T_52521 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,_T_52384}; // @[Mux.scala 19:72:@25180.4]
  assign _T_52523 = _T_2700 ? _T_52521 : 16'h0; // @[Mux.scala 19:72:@25181.4]
  assign _T_52538 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,_T_52401}; // @[Mux.scala 19:72:@25196.4]
  assign _T_52540 = _T_2701 ? _T_52538 : 16'h0; // @[Mux.scala 19:72:@25197.4]
  assign _T_52555 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,_T_52418}; // @[Mux.scala 19:72:@25212.4]
  assign _T_52557 = _T_2702 ? _T_52555 : 16'h0; // @[Mux.scala 19:72:@25213.4]
  assign _T_52572 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,_T_52435}; // @[Mux.scala 19:72:@25228.4]
  assign _T_52574 = _T_2703 ? _T_52572 : 16'h0; // @[Mux.scala 19:72:@25229.4]
  assign _T_52589 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,_T_52452}; // @[Mux.scala 19:72:@25244.4]
  assign _T_52591 = _T_2704 ? _T_52589 : 16'h0; // @[Mux.scala 19:72:@25245.4]
  assign _T_52592 = _T_52336 | _T_52353; // @[Mux.scala 19:72:@25246.4]
  assign _T_52593 = _T_52592 | _T_52370; // @[Mux.scala 19:72:@25247.4]
  assign _T_52594 = _T_52593 | _T_52387; // @[Mux.scala 19:72:@25248.4]
  assign _T_52595 = _T_52594 | _T_52404; // @[Mux.scala 19:72:@25249.4]
  assign _T_52596 = _T_52595 | _T_52421; // @[Mux.scala 19:72:@25250.4]
  assign _T_52597 = _T_52596 | _T_52438; // @[Mux.scala 19:72:@25251.4]
  assign _T_52598 = _T_52597 | _T_52455; // @[Mux.scala 19:72:@25252.4]
  assign _T_52599 = _T_52598 | _T_52472; // @[Mux.scala 19:72:@25253.4]
  assign _T_52600 = _T_52599 | _T_52489; // @[Mux.scala 19:72:@25254.4]
  assign _T_52601 = _T_52600 | _T_52506; // @[Mux.scala 19:72:@25255.4]
  assign _T_52602 = _T_52601 | _T_52523; // @[Mux.scala 19:72:@25256.4]
  assign _T_52603 = _T_52602 | _T_52540; // @[Mux.scala 19:72:@25257.4]
  assign _T_52604 = _T_52603 | _T_52557; // @[Mux.scala 19:72:@25258.4]
  assign _T_52605 = _T_52604 | _T_52574; // @[Mux.scala 19:72:@25259.4]
  assign _T_52606 = _T_52605 | _T_52591; // @[Mux.scala 19:72:@25260.4]
  assign _T_53184 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@25610.4]
  assign _T_53191 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8}; // @[Mux.scala 19:72:@25617.4]
  assign _T_53192 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,_T_53184}; // @[Mux.scala 19:72:@25618.4]
  assign _T_53194 = _T_2689 ? _T_53192 : 16'h0; // @[Mux.scala 19:72:@25619.4]
  assign _T_53201 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@25626.4]
  assign _T_53208 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9}; // @[Mux.scala 19:72:@25633.4]
  assign _T_53209 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,_T_53201}; // @[Mux.scala 19:72:@25634.4]
  assign _T_53211 = _T_2690 ? _T_53209 : 16'h0; // @[Mux.scala 19:72:@25635.4]
  assign _T_53218 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@25642.4]
  assign _T_53225 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10}; // @[Mux.scala 19:72:@25649.4]
  assign _T_53226 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,_T_53218}; // @[Mux.scala 19:72:@25650.4]
  assign _T_53228 = _T_2691 ? _T_53226 : 16'h0; // @[Mux.scala 19:72:@25651.4]
  assign _T_53235 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@25658.4]
  assign _T_53242 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11}; // @[Mux.scala 19:72:@25665.4]
  assign _T_53243 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,_T_53235}; // @[Mux.scala 19:72:@25666.4]
  assign _T_53245 = _T_2692 ? _T_53243 : 16'h0; // @[Mux.scala 19:72:@25667.4]
  assign _T_53252 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@25674.4]
  assign _T_53259 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12}; // @[Mux.scala 19:72:@25681.4]
  assign _T_53260 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,_T_53252}; // @[Mux.scala 19:72:@25682.4]
  assign _T_53262 = _T_2693 ? _T_53260 : 16'h0; // @[Mux.scala 19:72:@25683.4]
  assign _T_53269 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@25690.4]
  assign _T_53276 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13}; // @[Mux.scala 19:72:@25697.4]
  assign _T_53277 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,_T_53269}; // @[Mux.scala 19:72:@25698.4]
  assign _T_53279 = _T_2694 ? _T_53277 : 16'h0; // @[Mux.scala 19:72:@25699.4]
  assign _T_53286 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@25706.4]
  assign _T_53293 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14}; // @[Mux.scala 19:72:@25713.4]
  assign _T_53294 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,_T_53286}; // @[Mux.scala 19:72:@25714.4]
  assign _T_53296 = _T_2695 ? _T_53294 : 16'h0; // @[Mux.scala 19:72:@25715.4]
  assign _T_53303 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@25722.4]
  assign _T_53310 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15}; // @[Mux.scala 19:72:@25729.4]
  assign _T_53311 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,_T_53303}; // @[Mux.scala 19:72:@25730.4]
  assign _T_53313 = _T_2696 ? _T_53311 : 16'h0; // @[Mux.scala 19:72:@25731.4]
  assign _T_53328 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,_T_53191}; // @[Mux.scala 19:72:@25746.4]
  assign _T_53330 = _T_2697 ? _T_53328 : 16'h0; // @[Mux.scala 19:72:@25747.4]
  assign _T_53345 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,_T_53208}; // @[Mux.scala 19:72:@25762.4]
  assign _T_53347 = _T_2698 ? _T_53345 : 16'h0; // @[Mux.scala 19:72:@25763.4]
  assign _T_53362 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,_T_53225}; // @[Mux.scala 19:72:@25778.4]
  assign _T_53364 = _T_2699 ? _T_53362 : 16'h0; // @[Mux.scala 19:72:@25779.4]
  assign _T_53379 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,_T_53242}; // @[Mux.scala 19:72:@25794.4]
  assign _T_53381 = _T_2700 ? _T_53379 : 16'h0; // @[Mux.scala 19:72:@25795.4]
  assign _T_53396 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,_T_53259}; // @[Mux.scala 19:72:@25810.4]
  assign _T_53398 = _T_2701 ? _T_53396 : 16'h0; // @[Mux.scala 19:72:@25811.4]
  assign _T_53413 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,_T_53276}; // @[Mux.scala 19:72:@25826.4]
  assign _T_53415 = _T_2702 ? _T_53413 : 16'h0; // @[Mux.scala 19:72:@25827.4]
  assign _T_53430 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,_T_53293}; // @[Mux.scala 19:72:@25842.4]
  assign _T_53432 = _T_2703 ? _T_53430 : 16'h0; // @[Mux.scala 19:72:@25843.4]
  assign _T_53447 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,_T_53310}; // @[Mux.scala 19:72:@25858.4]
  assign _T_53449 = _T_2704 ? _T_53447 : 16'h0; // @[Mux.scala 19:72:@25859.4]
  assign _T_53450 = _T_53194 | _T_53211; // @[Mux.scala 19:72:@25860.4]
  assign _T_53451 = _T_53450 | _T_53228; // @[Mux.scala 19:72:@25861.4]
  assign _T_53452 = _T_53451 | _T_53245; // @[Mux.scala 19:72:@25862.4]
  assign _T_53453 = _T_53452 | _T_53262; // @[Mux.scala 19:72:@25863.4]
  assign _T_53454 = _T_53453 | _T_53279; // @[Mux.scala 19:72:@25864.4]
  assign _T_53455 = _T_53454 | _T_53296; // @[Mux.scala 19:72:@25865.4]
  assign _T_53456 = _T_53455 | _T_53313; // @[Mux.scala 19:72:@25866.4]
  assign _T_53457 = _T_53456 | _T_53330; // @[Mux.scala 19:72:@25867.4]
  assign _T_53458 = _T_53457 | _T_53347; // @[Mux.scala 19:72:@25868.4]
  assign _T_53459 = _T_53458 | _T_53364; // @[Mux.scala 19:72:@25869.4]
  assign _T_53460 = _T_53459 | _T_53381; // @[Mux.scala 19:72:@25870.4]
  assign _T_53461 = _T_53460 | _T_53398; // @[Mux.scala 19:72:@25871.4]
  assign _T_53462 = _T_53461 | _T_53415; // @[Mux.scala 19:72:@25872.4]
  assign _T_53463 = _T_53462 | _T_53432; // @[Mux.scala 19:72:@25873.4]
  assign _T_53464 = _T_53463 | _T_53449; // @[Mux.scala 19:72:@25874.4]
  assign _T_54042 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@26224.4]
  assign _T_54049 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8}; // @[Mux.scala 19:72:@26231.4]
  assign _T_54050 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,_T_54042}; // @[Mux.scala 19:72:@26232.4]
  assign _T_54052 = _T_2689 ? _T_54050 : 16'h0; // @[Mux.scala 19:72:@26233.4]
  assign _T_54059 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@26240.4]
  assign _T_54066 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9}; // @[Mux.scala 19:72:@26247.4]
  assign _T_54067 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,_T_54059}; // @[Mux.scala 19:72:@26248.4]
  assign _T_54069 = _T_2690 ? _T_54067 : 16'h0; // @[Mux.scala 19:72:@26249.4]
  assign _T_54076 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@26256.4]
  assign _T_54083 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10}; // @[Mux.scala 19:72:@26263.4]
  assign _T_54084 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,_T_54076}; // @[Mux.scala 19:72:@26264.4]
  assign _T_54086 = _T_2691 ? _T_54084 : 16'h0; // @[Mux.scala 19:72:@26265.4]
  assign _T_54093 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@26272.4]
  assign _T_54100 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11}; // @[Mux.scala 19:72:@26279.4]
  assign _T_54101 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,_T_54093}; // @[Mux.scala 19:72:@26280.4]
  assign _T_54103 = _T_2692 ? _T_54101 : 16'h0; // @[Mux.scala 19:72:@26281.4]
  assign _T_54110 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@26288.4]
  assign _T_54117 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12}; // @[Mux.scala 19:72:@26295.4]
  assign _T_54118 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,_T_54110}; // @[Mux.scala 19:72:@26296.4]
  assign _T_54120 = _T_2693 ? _T_54118 : 16'h0; // @[Mux.scala 19:72:@26297.4]
  assign _T_54127 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@26304.4]
  assign _T_54134 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13}; // @[Mux.scala 19:72:@26311.4]
  assign _T_54135 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,_T_54127}; // @[Mux.scala 19:72:@26312.4]
  assign _T_54137 = _T_2694 ? _T_54135 : 16'h0; // @[Mux.scala 19:72:@26313.4]
  assign _T_54144 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@26320.4]
  assign _T_54151 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14}; // @[Mux.scala 19:72:@26327.4]
  assign _T_54152 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,_T_54144}; // @[Mux.scala 19:72:@26328.4]
  assign _T_54154 = _T_2695 ? _T_54152 : 16'h0; // @[Mux.scala 19:72:@26329.4]
  assign _T_54161 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@26336.4]
  assign _T_54168 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15}; // @[Mux.scala 19:72:@26343.4]
  assign _T_54169 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,_T_54161}; // @[Mux.scala 19:72:@26344.4]
  assign _T_54171 = _T_2696 ? _T_54169 : 16'h0; // @[Mux.scala 19:72:@26345.4]
  assign _T_54186 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,_T_54049}; // @[Mux.scala 19:72:@26360.4]
  assign _T_54188 = _T_2697 ? _T_54186 : 16'h0; // @[Mux.scala 19:72:@26361.4]
  assign _T_54203 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,_T_54066}; // @[Mux.scala 19:72:@26376.4]
  assign _T_54205 = _T_2698 ? _T_54203 : 16'h0; // @[Mux.scala 19:72:@26377.4]
  assign _T_54220 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,_T_54083}; // @[Mux.scala 19:72:@26392.4]
  assign _T_54222 = _T_2699 ? _T_54220 : 16'h0; // @[Mux.scala 19:72:@26393.4]
  assign _T_54237 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,_T_54100}; // @[Mux.scala 19:72:@26408.4]
  assign _T_54239 = _T_2700 ? _T_54237 : 16'h0; // @[Mux.scala 19:72:@26409.4]
  assign _T_54254 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,_T_54117}; // @[Mux.scala 19:72:@26424.4]
  assign _T_54256 = _T_2701 ? _T_54254 : 16'h0; // @[Mux.scala 19:72:@26425.4]
  assign _T_54271 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,_T_54134}; // @[Mux.scala 19:72:@26440.4]
  assign _T_54273 = _T_2702 ? _T_54271 : 16'h0; // @[Mux.scala 19:72:@26441.4]
  assign _T_54288 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,_T_54151}; // @[Mux.scala 19:72:@26456.4]
  assign _T_54290 = _T_2703 ? _T_54288 : 16'h0; // @[Mux.scala 19:72:@26457.4]
  assign _T_54305 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,_T_54168}; // @[Mux.scala 19:72:@26472.4]
  assign _T_54307 = _T_2704 ? _T_54305 : 16'h0; // @[Mux.scala 19:72:@26473.4]
  assign _T_54308 = _T_54052 | _T_54069; // @[Mux.scala 19:72:@26474.4]
  assign _T_54309 = _T_54308 | _T_54086; // @[Mux.scala 19:72:@26475.4]
  assign _T_54310 = _T_54309 | _T_54103; // @[Mux.scala 19:72:@26476.4]
  assign _T_54311 = _T_54310 | _T_54120; // @[Mux.scala 19:72:@26477.4]
  assign _T_54312 = _T_54311 | _T_54137; // @[Mux.scala 19:72:@26478.4]
  assign _T_54313 = _T_54312 | _T_54154; // @[Mux.scala 19:72:@26479.4]
  assign _T_54314 = _T_54313 | _T_54171; // @[Mux.scala 19:72:@26480.4]
  assign _T_54315 = _T_54314 | _T_54188; // @[Mux.scala 19:72:@26481.4]
  assign _T_54316 = _T_54315 | _T_54205; // @[Mux.scala 19:72:@26482.4]
  assign _T_54317 = _T_54316 | _T_54222; // @[Mux.scala 19:72:@26483.4]
  assign _T_54318 = _T_54317 | _T_54239; // @[Mux.scala 19:72:@26484.4]
  assign _T_54319 = _T_54318 | _T_54256; // @[Mux.scala 19:72:@26485.4]
  assign _T_54320 = _T_54319 | _T_54273; // @[Mux.scala 19:72:@26486.4]
  assign _T_54321 = _T_54320 | _T_54290; // @[Mux.scala 19:72:@26487.4]
  assign _T_54322 = _T_54321 | _T_54307; // @[Mux.scala 19:72:@26488.4]
  assign _T_54900 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@26838.4]
  assign _T_54907 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8}; // @[Mux.scala 19:72:@26845.4]
  assign _T_54908 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,_T_54900}; // @[Mux.scala 19:72:@26846.4]
  assign _T_54910 = _T_2689 ? _T_54908 : 16'h0; // @[Mux.scala 19:72:@26847.4]
  assign _T_54917 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@26854.4]
  assign _T_54924 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9}; // @[Mux.scala 19:72:@26861.4]
  assign _T_54925 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,_T_54917}; // @[Mux.scala 19:72:@26862.4]
  assign _T_54927 = _T_2690 ? _T_54925 : 16'h0; // @[Mux.scala 19:72:@26863.4]
  assign _T_54934 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@26870.4]
  assign _T_54941 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10}; // @[Mux.scala 19:72:@26877.4]
  assign _T_54942 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,_T_54934}; // @[Mux.scala 19:72:@26878.4]
  assign _T_54944 = _T_2691 ? _T_54942 : 16'h0; // @[Mux.scala 19:72:@26879.4]
  assign _T_54951 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@26886.4]
  assign _T_54958 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11}; // @[Mux.scala 19:72:@26893.4]
  assign _T_54959 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,_T_54951}; // @[Mux.scala 19:72:@26894.4]
  assign _T_54961 = _T_2692 ? _T_54959 : 16'h0; // @[Mux.scala 19:72:@26895.4]
  assign _T_54968 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@26902.4]
  assign _T_54975 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12}; // @[Mux.scala 19:72:@26909.4]
  assign _T_54976 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,_T_54968}; // @[Mux.scala 19:72:@26910.4]
  assign _T_54978 = _T_2693 ? _T_54976 : 16'h0; // @[Mux.scala 19:72:@26911.4]
  assign _T_54985 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@26918.4]
  assign _T_54992 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13}; // @[Mux.scala 19:72:@26925.4]
  assign _T_54993 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,_T_54985}; // @[Mux.scala 19:72:@26926.4]
  assign _T_54995 = _T_2694 ? _T_54993 : 16'h0; // @[Mux.scala 19:72:@26927.4]
  assign _T_55002 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@26934.4]
  assign _T_55009 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14}; // @[Mux.scala 19:72:@26941.4]
  assign _T_55010 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,_T_55002}; // @[Mux.scala 19:72:@26942.4]
  assign _T_55012 = _T_2695 ? _T_55010 : 16'h0; // @[Mux.scala 19:72:@26943.4]
  assign _T_55019 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@26950.4]
  assign _T_55026 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15}; // @[Mux.scala 19:72:@26957.4]
  assign _T_55027 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,_T_55019}; // @[Mux.scala 19:72:@26958.4]
  assign _T_55029 = _T_2696 ? _T_55027 : 16'h0; // @[Mux.scala 19:72:@26959.4]
  assign _T_55044 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,_T_54907}; // @[Mux.scala 19:72:@26974.4]
  assign _T_55046 = _T_2697 ? _T_55044 : 16'h0; // @[Mux.scala 19:72:@26975.4]
  assign _T_55061 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,_T_54924}; // @[Mux.scala 19:72:@26990.4]
  assign _T_55063 = _T_2698 ? _T_55061 : 16'h0; // @[Mux.scala 19:72:@26991.4]
  assign _T_55078 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,_T_54941}; // @[Mux.scala 19:72:@27006.4]
  assign _T_55080 = _T_2699 ? _T_55078 : 16'h0; // @[Mux.scala 19:72:@27007.4]
  assign _T_55095 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,_T_54958}; // @[Mux.scala 19:72:@27022.4]
  assign _T_55097 = _T_2700 ? _T_55095 : 16'h0; // @[Mux.scala 19:72:@27023.4]
  assign _T_55112 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,_T_54975}; // @[Mux.scala 19:72:@27038.4]
  assign _T_55114 = _T_2701 ? _T_55112 : 16'h0; // @[Mux.scala 19:72:@27039.4]
  assign _T_55129 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,_T_54992}; // @[Mux.scala 19:72:@27054.4]
  assign _T_55131 = _T_2702 ? _T_55129 : 16'h0; // @[Mux.scala 19:72:@27055.4]
  assign _T_55146 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,_T_55009}; // @[Mux.scala 19:72:@27070.4]
  assign _T_55148 = _T_2703 ? _T_55146 : 16'h0; // @[Mux.scala 19:72:@27071.4]
  assign _T_55163 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,_T_55026}; // @[Mux.scala 19:72:@27086.4]
  assign _T_55165 = _T_2704 ? _T_55163 : 16'h0; // @[Mux.scala 19:72:@27087.4]
  assign _T_55166 = _T_54910 | _T_54927; // @[Mux.scala 19:72:@27088.4]
  assign _T_55167 = _T_55166 | _T_54944; // @[Mux.scala 19:72:@27089.4]
  assign _T_55168 = _T_55167 | _T_54961; // @[Mux.scala 19:72:@27090.4]
  assign _T_55169 = _T_55168 | _T_54978; // @[Mux.scala 19:72:@27091.4]
  assign _T_55170 = _T_55169 | _T_54995; // @[Mux.scala 19:72:@27092.4]
  assign _T_55171 = _T_55170 | _T_55012; // @[Mux.scala 19:72:@27093.4]
  assign _T_55172 = _T_55171 | _T_55029; // @[Mux.scala 19:72:@27094.4]
  assign _T_55173 = _T_55172 | _T_55046; // @[Mux.scala 19:72:@27095.4]
  assign _T_55174 = _T_55173 | _T_55063; // @[Mux.scala 19:72:@27096.4]
  assign _T_55175 = _T_55174 | _T_55080; // @[Mux.scala 19:72:@27097.4]
  assign _T_55176 = _T_55175 | _T_55097; // @[Mux.scala 19:72:@27098.4]
  assign _T_55177 = _T_55176 | _T_55114; // @[Mux.scala 19:72:@27099.4]
  assign _T_55178 = _T_55177 | _T_55131; // @[Mux.scala 19:72:@27100.4]
  assign _T_55179 = _T_55178 | _T_55148; // @[Mux.scala 19:72:@27101.4]
  assign _T_55180 = _T_55179 | _T_55165; // @[Mux.scala 19:72:@27102.4]
  assign _T_55758 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@27452.4]
  assign _T_55765 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8}; // @[Mux.scala 19:72:@27459.4]
  assign _T_55766 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,_T_55758}; // @[Mux.scala 19:72:@27460.4]
  assign _T_55768 = _T_2689 ? _T_55766 : 16'h0; // @[Mux.scala 19:72:@27461.4]
  assign _T_55775 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@27468.4]
  assign _T_55782 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9}; // @[Mux.scala 19:72:@27475.4]
  assign _T_55783 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,_T_55775}; // @[Mux.scala 19:72:@27476.4]
  assign _T_55785 = _T_2690 ? _T_55783 : 16'h0; // @[Mux.scala 19:72:@27477.4]
  assign _T_55792 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@27484.4]
  assign _T_55799 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10}; // @[Mux.scala 19:72:@27491.4]
  assign _T_55800 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,_T_55792}; // @[Mux.scala 19:72:@27492.4]
  assign _T_55802 = _T_2691 ? _T_55800 : 16'h0; // @[Mux.scala 19:72:@27493.4]
  assign _T_55809 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@27500.4]
  assign _T_55816 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11}; // @[Mux.scala 19:72:@27507.4]
  assign _T_55817 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,_T_55809}; // @[Mux.scala 19:72:@27508.4]
  assign _T_55819 = _T_2692 ? _T_55817 : 16'h0; // @[Mux.scala 19:72:@27509.4]
  assign _T_55826 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@27516.4]
  assign _T_55833 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12}; // @[Mux.scala 19:72:@27523.4]
  assign _T_55834 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,_T_55826}; // @[Mux.scala 19:72:@27524.4]
  assign _T_55836 = _T_2693 ? _T_55834 : 16'h0; // @[Mux.scala 19:72:@27525.4]
  assign _T_55843 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@27532.4]
  assign _T_55850 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13}; // @[Mux.scala 19:72:@27539.4]
  assign _T_55851 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,_T_55843}; // @[Mux.scala 19:72:@27540.4]
  assign _T_55853 = _T_2694 ? _T_55851 : 16'h0; // @[Mux.scala 19:72:@27541.4]
  assign _T_55860 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@27548.4]
  assign _T_55867 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14}; // @[Mux.scala 19:72:@27555.4]
  assign _T_55868 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,_T_55860}; // @[Mux.scala 19:72:@27556.4]
  assign _T_55870 = _T_2695 ? _T_55868 : 16'h0; // @[Mux.scala 19:72:@27557.4]
  assign _T_55877 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@27564.4]
  assign _T_55884 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15}; // @[Mux.scala 19:72:@27571.4]
  assign _T_55885 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,_T_55877}; // @[Mux.scala 19:72:@27572.4]
  assign _T_55887 = _T_2696 ? _T_55885 : 16'h0; // @[Mux.scala 19:72:@27573.4]
  assign _T_55902 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,_T_55765}; // @[Mux.scala 19:72:@27588.4]
  assign _T_55904 = _T_2697 ? _T_55902 : 16'h0; // @[Mux.scala 19:72:@27589.4]
  assign _T_55919 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,_T_55782}; // @[Mux.scala 19:72:@27604.4]
  assign _T_55921 = _T_2698 ? _T_55919 : 16'h0; // @[Mux.scala 19:72:@27605.4]
  assign _T_55936 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,_T_55799}; // @[Mux.scala 19:72:@27620.4]
  assign _T_55938 = _T_2699 ? _T_55936 : 16'h0; // @[Mux.scala 19:72:@27621.4]
  assign _T_55953 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,_T_55816}; // @[Mux.scala 19:72:@27636.4]
  assign _T_55955 = _T_2700 ? _T_55953 : 16'h0; // @[Mux.scala 19:72:@27637.4]
  assign _T_55970 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,_T_55833}; // @[Mux.scala 19:72:@27652.4]
  assign _T_55972 = _T_2701 ? _T_55970 : 16'h0; // @[Mux.scala 19:72:@27653.4]
  assign _T_55987 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,_T_55850}; // @[Mux.scala 19:72:@27668.4]
  assign _T_55989 = _T_2702 ? _T_55987 : 16'h0; // @[Mux.scala 19:72:@27669.4]
  assign _T_56004 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,_T_55867}; // @[Mux.scala 19:72:@27684.4]
  assign _T_56006 = _T_2703 ? _T_56004 : 16'h0; // @[Mux.scala 19:72:@27685.4]
  assign _T_56021 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,_T_55884}; // @[Mux.scala 19:72:@27700.4]
  assign _T_56023 = _T_2704 ? _T_56021 : 16'h0; // @[Mux.scala 19:72:@27701.4]
  assign _T_56024 = _T_55768 | _T_55785; // @[Mux.scala 19:72:@27702.4]
  assign _T_56025 = _T_56024 | _T_55802; // @[Mux.scala 19:72:@27703.4]
  assign _T_56026 = _T_56025 | _T_55819; // @[Mux.scala 19:72:@27704.4]
  assign _T_56027 = _T_56026 | _T_55836; // @[Mux.scala 19:72:@27705.4]
  assign _T_56028 = _T_56027 | _T_55853; // @[Mux.scala 19:72:@27706.4]
  assign _T_56029 = _T_56028 | _T_55870; // @[Mux.scala 19:72:@27707.4]
  assign _T_56030 = _T_56029 | _T_55887; // @[Mux.scala 19:72:@27708.4]
  assign _T_56031 = _T_56030 | _T_55904; // @[Mux.scala 19:72:@27709.4]
  assign _T_56032 = _T_56031 | _T_55921; // @[Mux.scala 19:72:@27710.4]
  assign _T_56033 = _T_56032 | _T_55938; // @[Mux.scala 19:72:@27711.4]
  assign _T_56034 = _T_56033 | _T_55955; // @[Mux.scala 19:72:@27712.4]
  assign _T_56035 = _T_56034 | _T_55972; // @[Mux.scala 19:72:@27713.4]
  assign _T_56036 = _T_56035 | _T_55989; // @[Mux.scala 19:72:@27714.4]
  assign _T_56037 = _T_56036 | _T_56006; // @[Mux.scala 19:72:@27715.4]
  assign _T_56038 = _T_56037 | _T_56023; // @[Mux.scala 19:72:@27716.4]
  assign _T_56616 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@28066.4]
  assign _T_56623 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8}; // @[Mux.scala 19:72:@28073.4]
  assign _T_56624 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,_T_56616}; // @[Mux.scala 19:72:@28074.4]
  assign _T_56626 = _T_2689 ? _T_56624 : 16'h0; // @[Mux.scala 19:72:@28075.4]
  assign _T_56633 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@28082.4]
  assign _T_56640 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9}; // @[Mux.scala 19:72:@28089.4]
  assign _T_56641 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,_T_56633}; // @[Mux.scala 19:72:@28090.4]
  assign _T_56643 = _T_2690 ? _T_56641 : 16'h0; // @[Mux.scala 19:72:@28091.4]
  assign _T_56650 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@28098.4]
  assign _T_56657 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10}; // @[Mux.scala 19:72:@28105.4]
  assign _T_56658 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,_T_56650}; // @[Mux.scala 19:72:@28106.4]
  assign _T_56660 = _T_2691 ? _T_56658 : 16'h0; // @[Mux.scala 19:72:@28107.4]
  assign _T_56667 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@28114.4]
  assign _T_56674 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11}; // @[Mux.scala 19:72:@28121.4]
  assign _T_56675 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,_T_56667}; // @[Mux.scala 19:72:@28122.4]
  assign _T_56677 = _T_2692 ? _T_56675 : 16'h0; // @[Mux.scala 19:72:@28123.4]
  assign _T_56684 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@28130.4]
  assign _T_56691 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12}; // @[Mux.scala 19:72:@28137.4]
  assign _T_56692 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,_T_56684}; // @[Mux.scala 19:72:@28138.4]
  assign _T_56694 = _T_2693 ? _T_56692 : 16'h0; // @[Mux.scala 19:72:@28139.4]
  assign _T_56701 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@28146.4]
  assign _T_56708 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13}; // @[Mux.scala 19:72:@28153.4]
  assign _T_56709 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,_T_56701}; // @[Mux.scala 19:72:@28154.4]
  assign _T_56711 = _T_2694 ? _T_56709 : 16'h0; // @[Mux.scala 19:72:@28155.4]
  assign _T_56718 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@28162.4]
  assign _T_56725 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14}; // @[Mux.scala 19:72:@28169.4]
  assign _T_56726 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,_T_56718}; // @[Mux.scala 19:72:@28170.4]
  assign _T_56728 = _T_2695 ? _T_56726 : 16'h0; // @[Mux.scala 19:72:@28171.4]
  assign _T_56735 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@28178.4]
  assign _T_56742 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15}; // @[Mux.scala 19:72:@28185.4]
  assign _T_56743 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,_T_56735}; // @[Mux.scala 19:72:@28186.4]
  assign _T_56745 = _T_2696 ? _T_56743 : 16'h0; // @[Mux.scala 19:72:@28187.4]
  assign _T_56760 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,_T_56623}; // @[Mux.scala 19:72:@28202.4]
  assign _T_56762 = _T_2697 ? _T_56760 : 16'h0; // @[Mux.scala 19:72:@28203.4]
  assign _T_56777 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,_T_56640}; // @[Mux.scala 19:72:@28218.4]
  assign _T_56779 = _T_2698 ? _T_56777 : 16'h0; // @[Mux.scala 19:72:@28219.4]
  assign _T_56794 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,_T_56657}; // @[Mux.scala 19:72:@28234.4]
  assign _T_56796 = _T_2699 ? _T_56794 : 16'h0; // @[Mux.scala 19:72:@28235.4]
  assign _T_56811 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,_T_56674}; // @[Mux.scala 19:72:@28250.4]
  assign _T_56813 = _T_2700 ? _T_56811 : 16'h0; // @[Mux.scala 19:72:@28251.4]
  assign _T_56828 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,_T_56691}; // @[Mux.scala 19:72:@28266.4]
  assign _T_56830 = _T_2701 ? _T_56828 : 16'h0; // @[Mux.scala 19:72:@28267.4]
  assign _T_56845 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,_T_56708}; // @[Mux.scala 19:72:@28282.4]
  assign _T_56847 = _T_2702 ? _T_56845 : 16'h0; // @[Mux.scala 19:72:@28283.4]
  assign _T_56862 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,_T_56725}; // @[Mux.scala 19:72:@28298.4]
  assign _T_56864 = _T_2703 ? _T_56862 : 16'h0; // @[Mux.scala 19:72:@28299.4]
  assign _T_56879 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,_T_56742}; // @[Mux.scala 19:72:@28314.4]
  assign _T_56881 = _T_2704 ? _T_56879 : 16'h0; // @[Mux.scala 19:72:@28315.4]
  assign _T_56882 = _T_56626 | _T_56643; // @[Mux.scala 19:72:@28316.4]
  assign _T_56883 = _T_56882 | _T_56660; // @[Mux.scala 19:72:@28317.4]
  assign _T_56884 = _T_56883 | _T_56677; // @[Mux.scala 19:72:@28318.4]
  assign _T_56885 = _T_56884 | _T_56694; // @[Mux.scala 19:72:@28319.4]
  assign _T_56886 = _T_56885 | _T_56711; // @[Mux.scala 19:72:@28320.4]
  assign _T_56887 = _T_56886 | _T_56728; // @[Mux.scala 19:72:@28321.4]
  assign _T_56888 = _T_56887 | _T_56745; // @[Mux.scala 19:72:@28322.4]
  assign _T_56889 = _T_56888 | _T_56762; // @[Mux.scala 19:72:@28323.4]
  assign _T_56890 = _T_56889 | _T_56779; // @[Mux.scala 19:72:@28324.4]
  assign _T_56891 = _T_56890 | _T_56796; // @[Mux.scala 19:72:@28325.4]
  assign _T_56892 = _T_56891 | _T_56813; // @[Mux.scala 19:72:@28326.4]
  assign _T_56893 = _T_56892 | _T_56830; // @[Mux.scala 19:72:@28327.4]
  assign _T_56894 = _T_56893 | _T_56847; // @[Mux.scala 19:72:@28328.4]
  assign _T_56895 = _T_56894 | _T_56864; // @[Mux.scala 19:72:@28329.4]
  assign _T_56896 = _T_56895 | _T_56881; // @[Mux.scala 19:72:@28330.4]
  assign _T_57474 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@28680.4]
  assign _T_57481 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8}; // @[Mux.scala 19:72:@28687.4]
  assign _T_57482 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,_T_57474}; // @[Mux.scala 19:72:@28688.4]
  assign _T_57484 = _T_2689 ? _T_57482 : 16'h0; // @[Mux.scala 19:72:@28689.4]
  assign _T_57491 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@28696.4]
  assign _T_57498 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9}; // @[Mux.scala 19:72:@28703.4]
  assign _T_57499 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,_T_57491}; // @[Mux.scala 19:72:@28704.4]
  assign _T_57501 = _T_2690 ? _T_57499 : 16'h0; // @[Mux.scala 19:72:@28705.4]
  assign _T_57508 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@28712.4]
  assign _T_57515 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10}; // @[Mux.scala 19:72:@28719.4]
  assign _T_57516 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,_T_57508}; // @[Mux.scala 19:72:@28720.4]
  assign _T_57518 = _T_2691 ? _T_57516 : 16'h0; // @[Mux.scala 19:72:@28721.4]
  assign _T_57525 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@28728.4]
  assign _T_57532 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11}; // @[Mux.scala 19:72:@28735.4]
  assign _T_57533 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,_T_57525}; // @[Mux.scala 19:72:@28736.4]
  assign _T_57535 = _T_2692 ? _T_57533 : 16'h0; // @[Mux.scala 19:72:@28737.4]
  assign _T_57542 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@28744.4]
  assign _T_57549 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12}; // @[Mux.scala 19:72:@28751.4]
  assign _T_57550 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,_T_57542}; // @[Mux.scala 19:72:@28752.4]
  assign _T_57552 = _T_2693 ? _T_57550 : 16'h0; // @[Mux.scala 19:72:@28753.4]
  assign _T_57559 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@28760.4]
  assign _T_57566 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13}; // @[Mux.scala 19:72:@28767.4]
  assign _T_57567 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,_T_57559}; // @[Mux.scala 19:72:@28768.4]
  assign _T_57569 = _T_2694 ? _T_57567 : 16'h0; // @[Mux.scala 19:72:@28769.4]
  assign _T_57576 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@28776.4]
  assign _T_57583 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14}; // @[Mux.scala 19:72:@28783.4]
  assign _T_57584 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,_T_57576}; // @[Mux.scala 19:72:@28784.4]
  assign _T_57586 = _T_2695 ? _T_57584 : 16'h0; // @[Mux.scala 19:72:@28785.4]
  assign _T_57593 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@28792.4]
  assign _T_57600 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15}; // @[Mux.scala 19:72:@28799.4]
  assign _T_57601 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,_T_57593}; // @[Mux.scala 19:72:@28800.4]
  assign _T_57603 = _T_2696 ? _T_57601 : 16'h0; // @[Mux.scala 19:72:@28801.4]
  assign _T_57618 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,_T_57481}; // @[Mux.scala 19:72:@28816.4]
  assign _T_57620 = _T_2697 ? _T_57618 : 16'h0; // @[Mux.scala 19:72:@28817.4]
  assign _T_57635 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,_T_57498}; // @[Mux.scala 19:72:@28832.4]
  assign _T_57637 = _T_2698 ? _T_57635 : 16'h0; // @[Mux.scala 19:72:@28833.4]
  assign _T_57652 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,_T_57515}; // @[Mux.scala 19:72:@28848.4]
  assign _T_57654 = _T_2699 ? _T_57652 : 16'h0; // @[Mux.scala 19:72:@28849.4]
  assign _T_57669 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,_T_57532}; // @[Mux.scala 19:72:@28864.4]
  assign _T_57671 = _T_2700 ? _T_57669 : 16'h0; // @[Mux.scala 19:72:@28865.4]
  assign _T_57686 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,_T_57549}; // @[Mux.scala 19:72:@28880.4]
  assign _T_57688 = _T_2701 ? _T_57686 : 16'h0; // @[Mux.scala 19:72:@28881.4]
  assign _T_57703 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,_T_57566}; // @[Mux.scala 19:72:@28896.4]
  assign _T_57705 = _T_2702 ? _T_57703 : 16'h0; // @[Mux.scala 19:72:@28897.4]
  assign _T_57720 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,_T_57583}; // @[Mux.scala 19:72:@28912.4]
  assign _T_57722 = _T_2703 ? _T_57720 : 16'h0; // @[Mux.scala 19:72:@28913.4]
  assign _T_57737 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,_T_57600}; // @[Mux.scala 19:72:@28928.4]
  assign _T_57739 = _T_2704 ? _T_57737 : 16'h0; // @[Mux.scala 19:72:@28929.4]
  assign _T_57740 = _T_57484 | _T_57501; // @[Mux.scala 19:72:@28930.4]
  assign _T_57741 = _T_57740 | _T_57518; // @[Mux.scala 19:72:@28931.4]
  assign _T_57742 = _T_57741 | _T_57535; // @[Mux.scala 19:72:@28932.4]
  assign _T_57743 = _T_57742 | _T_57552; // @[Mux.scala 19:72:@28933.4]
  assign _T_57744 = _T_57743 | _T_57569; // @[Mux.scala 19:72:@28934.4]
  assign _T_57745 = _T_57744 | _T_57586; // @[Mux.scala 19:72:@28935.4]
  assign _T_57746 = _T_57745 | _T_57603; // @[Mux.scala 19:72:@28936.4]
  assign _T_57747 = _T_57746 | _T_57620; // @[Mux.scala 19:72:@28937.4]
  assign _T_57748 = _T_57747 | _T_57637; // @[Mux.scala 19:72:@28938.4]
  assign _T_57749 = _T_57748 | _T_57654; // @[Mux.scala 19:72:@28939.4]
  assign _T_57750 = _T_57749 | _T_57671; // @[Mux.scala 19:72:@28940.4]
  assign _T_57751 = _T_57750 | _T_57688; // @[Mux.scala 19:72:@28941.4]
  assign _T_57752 = _T_57751 | _T_57705; // @[Mux.scala 19:72:@28942.4]
  assign _T_57753 = _T_57752 | _T_57722; // @[Mux.scala 19:72:@28943.4]
  assign _T_57754 = _T_57753 | _T_57739; // @[Mux.scala 19:72:@28944.4]
  assign _T_58332 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@29294.4]
  assign _T_58339 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8}; // @[Mux.scala 19:72:@29301.4]
  assign _T_58340 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,_T_58332}; // @[Mux.scala 19:72:@29302.4]
  assign _T_58342 = _T_2689 ? _T_58340 : 16'h0; // @[Mux.scala 19:72:@29303.4]
  assign _T_58349 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@29310.4]
  assign _T_58356 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9}; // @[Mux.scala 19:72:@29317.4]
  assign _T_58357 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,_T_58349}; // @[Mux.scala 19:72:@29318.4]
  assign _T_58359 = _T_2690 ? _T_58357 : 16'h0; // @[Mux.scala 19:72:@29319.4]
  assign _T_58366 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@29326.4]
  assign _T_58373 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10}; // @[Mux.scala 19:72:@29333.4]
  assign _T_58374 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,_T_58366}; // @[Mux.scala 19:72:@29334.4]
  assign _T_58376 = _T_2691 ? _T_58374 : 16'h0; // @[Mux.scala 19:72:@29335.4]
  assign _T_58383 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@29342.4]
  assign _T_58390 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11}; // @[Mux.scala 19:72:@29349.4]
  assign _T_58391 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,_T_58383}; // @[Mux.scala 19:72:@29350.4]
  assign _T_58393 = _T_2692 ? _T_58391 : 16'h0; // @[Mux.scala 19:72:@29351.4]
  assign _T_58400 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@29358.4]
  assign _T_58407 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12}; // @[Mux.scala 19:72:@29365.4]
  assign _T_58408 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,_T_58400}; // @[Mux.scala 19:72:@29366.4]
  assign _T_58410 = _T_2693 ? _T_58408 : 16'h0; // @[Mux.scala 19:72:@29367.4]
  assign _T_58417 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@29374.4]
  assign _T_58424 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13}; // @[Mux.scala 19:72:@29381.4]
  assign _T_58425 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,_T_58417}; // @[Mux.scala 19:72:@29382.4]
  assign _T_58427 = _T_2694 ? _T_58425 : 16'h0; // @[Mux.scala 19:72:@29383.4]
  assign _T_58434 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@29390.4]
  assign _T_58441 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14}; // @[Mux.scala 19:72:@29397.4]
  assign _T_58442 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,_T_58434}; // @[Mux.scala 19:72:@29398.4]
  assign _T_58444 = _T_2695 ? _T_58442 : 16'h0; // @[Mux.scala 19:72:@29399.4]
  assign _T_58451 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@29406.4]
  assign _T_58458 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15}; // @[Mux.scala 19:72:@29413.4]
  assign _T_58459 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,_T_58451}; // @[Mux.scala 19:72:@29414.4]
  assign _T_58461 = _T_2696 ? _T_58459 : 16'h0; // @[Mux.scala 19:72:@29415.4]
  assign _T_58476 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,_T_58339}; // @[Mux.scala 19:72:@29430.4]
  assign _T_58478 = _T_2697 ? _T_58476 : 16'h0; // @[Mux.scala 19:72:@29431.4]
  assign _T_58493 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,_T_58356}; // @[Mux.scala 19:72:@29446.4]
  assign _T_58495 = _T_2698 ? _T_58493 : 16'h0; // @[Mux.scala 19:72:@29447.4]
  assign _T_58510 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,_T_58373}; // @[Mux.scala 19:72:@29462.4]
  assign _T_58512 = _T_2699 ? _T_58510 : 16'h0; // @[Mux.scala 19:72:@29463.4]
  assign _T_58527 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,_T_58390}; // @[Mux.scala 19:72:@29478.4]
  assign _T_58529 = _T_2700 ? _T_58527 : 16'h0; // @[Mux.scala 19:72:@29479.4]
  assign _T_58544 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,_T_58407}; // @[Mux.scala 19:72:@29494.4]
  assign _T_58546 = _T_2701 ? _T_58544 : 16'h0; // @[Mux.scala 19:72:@29495.4]
  assign _T_58561 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,_T_58424}; // @[Mux.scala 19:72:@29510.4]
  assign _T_58563 = _T_2702 ? _T_58561 : 16'h0; // @[Mux.scala 19:72:@29511.4]
  assign _T_58578 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,_T_58441}; // @[Mux.scala 19:72:@29526.4]
  assign _T_58580 = _T_2703 ? _T_58578 : 16'h0; // @[Mux.scala 19:72:@29527.4]
  assign _T_58595 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,_T_58458}; // @[Mux.scala 19:72:@29542.4]
  assign _T_58597 = _T_2704 ? _T_58595 : 16'h0; // @[Mux.scala 19:72:@29543.4]
  assign _T_58598 = _T_58342 | _T_58359; // @[Mux.scala 19:72:@29544.4]
  assign _T_58599 = _T_58598 | _T_58376; // @[Mux.scala 19:72:@29545.4]
  assign _T_58600 = _T_58599 | _T_58393; // @[Mux.scala 19:72:@29546.4]
  assign _T_58601 = _T_58600 | _T_58410; // @[Mux.scala 19:72:@29547.4]
  assign _T_58602 = _T_58601 | _T_58427; // @[Mux.scala 19:72:@29548.4]
  assign _T_58603 = _T_58602 | _T_58444; // @[Mux.scala 19:72:@29549.4]
  assign _T_58604 = _T_58603 | _T_58461; // @[Mux.scala 19:72:@29550.4]
  assign _T_58605 = _T_58604 | _T_58478; // @[Mux.scala 19:72:@29551.4]
  assign _T_58606 = _T_58605 | _T_58495; // @[Mux.scala 19:72:@29552.4]
  assign _T_58607 = _T_58606 | _T_58512; // @[Mux.scala 19:72:@29553.4]
  assign _T_58608 = _T_58607 | _T_58529; // @[Mux.scala 19:72:@29554.4]
  assign _T_58609 = _T_58608 | _T_58546; // @[Mux.scala 19:72:@29555.4]
  assign _T_58610 = _T_58609 | _T_58563; // @[Mux.scala 19:72:@29556.4]
  assign _T_58611 = _T_58610 | _T_58580; // @[Mux.scala 19:72:@29557.4]
  assign _T_58612 = _T_58611 | _T_58597; // @[Mux.scala 19:72:@29558.4]
  assign _T_59190 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0}; // @[Mux.scala 19:72:@29908.4]
  assign _T_59197 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8}; // @[Mux.scala 19:72:@29915.4]
  assign _T_59198 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,_T_59190}; // @[Mux.scala 19:72:@29916.4]
  assign _T_59200 = _T_2689 ? _T_59198 : 16'h0; // @[Mux.scala 19:72:@29917.4]
  assign _T_59207 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1}; // @[Mux.scala 19:72:@29924.4]
  assign _T_59214 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9}; // @[Mux.scala 19:72:@29931.4]
  assign _T_59215 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,_T_59207}; // @[Mux.scala 19:72:@29932.4]
  assign _T_59217 = _T_2690 ? _T_59215 : 16'h0; // @[Mux.scala 19:72:@29933.4]
  assign _T_59224 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2}; // @[Mux.scala 19:72:@29940.4]
  assign _T_59231 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10}; // @[Mux.scala 19:72:@29947.4]
  assign _T_59232 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,_T_59224}; // @[Mux.scala 19:72:@29948.4]
  assign _T_59234 = _T_2691 ? _T_59232 : 16'h0; // @[Mux.scala 19:72:@29949.4]
  assign _T_59241 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3}; // @[Mux.scala 19:72:@29956.4]
  assign _T_59248 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11}; // @[Mux.scala 19:72:@29963.4]
  assign _T_59249 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,_T_59241}; // @[Mux.scala 19:72:@29964.4]
  assign _T_59251 = _T_2692 ? _T_59249 : 16'h0; // @[Mux.scala 19:72:@29965.4]
  assign _T_59258 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4}; // @[Mux.scala 19:72:@29972.4]
  assign _T_59265 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12}; // @[Mux.scala 19:72:@29979.4]
  assign _T_59266 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,_T_59258}; // @[Mux.scala 19:72:@29980.4]
  assign _T_59268 = _T_2693 ? _T_59266 : 16'h0; // @[Mux.scala 19:72:@29981.4]
  assign _T_59275 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5}; // @[Mux.scala 19:72:@29988.4]
  assign _T_59282 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13}; // @[Mux.scala 19:72:@29995.4]
  assign _T_59283 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,_T_59275}; // @[Mux.scala 19:72:@29996.4]
  assign _T_59285 = _T_2694 ? _T_59283 : 16'h0; // @[Mux.scala 19:72:@29997.4]
  assign _T_59292 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6}; // @[Mux.scala 19:72:@30004.4]
  assign _T_59299 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14}; // @[Mux.scala 19:72:@30011.4]
  assign _T_59300 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,_T_59292}; // @[Mux.scala 19:72:@30012.4]
  assign _T_59302 = _T_2695 ? _T_59300 : 16'h0; // @[Mux.scala 19:72:@30013.4]
  assign _T_59309 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7}; // @[Mux.scala 19:72:@30020.4]
  assign _T_59316 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15}; // @[Mux.scala 19:72:@30027.4]
  assign _T_59317 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,_T_59309}; // @[Mux.scala 19:72:@30028.4]
  assign _T_59319 = _T_2696 ? _T_59317 : 16'h0; // @[Mux.scala 19:72:@30029.4]
  assign _T_59334 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,_T_59197}; // @[Mux.scala 19:72:@30044.4]
  assign _T_59336 = _T_2697 ? _T_59334 : 16'h0; // @[Mux.scala 19:72:@30045.4]
  assign _T_59351 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,_T_59214}; // @[Mux.scala 19:72:@30060.4]
  assign _T_59353 = _T_2698 ? _T_59351 : 16'h0; // @[Mux.scala 19:72:@30061.4]
  assign _T_59368 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,_T_59231}; // @[Mux.scala 19:72:@30076.4]
  assign _T_59370 = _T_2699 ? _T_59368 : 16'h0; // @[Mux.scala 19:72:@30077.4]
  assign _T_59385 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,_T_59248}; // @[Mux.scala 19:72:@30092.4]
  assign _T_59387 = _T_2700 ? _T_59385 : 16'h0; // @[Mux.scala 19:72:@30093.4]
  assign _T_59402 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,_T_59265}; // @[Mux.scala 19:72:@30108.4]
  assign _T_59404 = _T_2701 ? _T_59402 : 16'h0; // @[Mux.scala 19:72:@30109.4]
  assign _T_59419 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,_T_59282}; // @[Mux.scala 19:72:@30124.4]
  assign _T_59421 = _T_2702 ? _T_59419 : 16'h0; // @[Mux.scala 19:72:@30125.4]
  assign _T_59436 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,_T_59299}; // @[Mux.scala 19:72:@30140.4]
  assign _T_59438 = _T_2703 ? _T_59436 : 16'h0; // @[Mux.scala 19:72:@30141.4]
  assign _T_59453 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,_T_59316}; // @[Mux.scala 19:72:@30156.4]
  assign _T_59455 = _T_2704 ? _T_59453 : 16'h0; // @[Mux.scala 19:72:@30157.4]
  assign _T_59456 = _T_59200 | _T_59217; // @[Mux.scala 19:72:@30158.4]
  assign _T_59457 = _T_59456 | _T_59234; // @[Mux.scala 19:72:@30159.4]
  assign _T_59458 = _T_59457 | _T_59251; // @[Mux.scala 19:72:@30160.4]
  assign _T_59459 = _T_59458 | _T_59268; // @[Mux.scala 19:72:@30161.4]
  assign _T_59460 = _T_59459 | _T_59285; // @[Mux.scala 19:72:@30162.4]
  assign _T_59461 = _T_59460 | _T_59302; // @[Mux.scala 19:72:@30163.4]
  assign _T_59462 = _T_59461 | _T_59319; // @[Mux.scala 19:72:@30164.4]
  assign _T_59463 = _T_59462 | _T_59336; // @[Mux.scala 19:72:@30165.4]
  assign _T_59464 = _T_59463 | _T_59353; // @[Mux.scala 19:72:@30166.4]
  assign _T_59465 = _T_59464 | _T_59370; // @[Mux.scala 19:72:@30167.4]
  assign _T_59466 = _T_59465 | _T_59387; // @[Mux.scala 19:72:@30168.4]
  assign _T_59467 = _T_59466 | _T_59404; // @[Mux.scala 19:72:@30169.4]
  assign _T_59468 = _T_59467 | _T_59421; // @[Mux.scala 19:72:@30170.4]
  assign _T_59469 = _T_59468 | _T_59438; // @[Mux.scala 19:72:@30171.4]
  assign _T_59470 = _T_59469 | _T_59455; // @[Mux.scala 19:72:@30172.4]
  assign _T_60048 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0}; // @[Mux.scala 19:72:@30522.4]
  assign _T_60055 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8}; // @[Mux.scala 19:72:@30529.4]
  assign _T_60056 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,_T_60048}; // @[Mux.scala 19:72:@30530.4]
  assign _T_60058 = _T_2689 ? _T_60056 : 16'h0; // @[Mux.scala 19:72:@30531.4]
  assign _T_60065 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1}; // @[Mux.scala 19:72:@30538.4]
  assign _T_60072 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9}; // @[Mux.scala 19:72:@30545.4]
  assign _T_60073 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,_T_60065}; // @[Mux.scala 19:72:@30546.4]
  assign _T_60075 = _T_2690 ? _T_60073 : 16'h0; // @[Mux.scala 19:72:@30547.4]
  assign _T_60082 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2}; // @[Mux.scala 19:72:@30554.4]
  assign _T_60089 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10}; // @[Mux.scala 19:72:@30561.4]
  assign _T_60090 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,_T_60082}; // @[Mux.scala 19:72:@30562.4]
  assign _T_60092 = _T_2691 ? _T_60090 : 16'h0; // @[Mux.scala 19:72:@30563.4]
  assign _T_60099 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3}; // @[Mux.scala 19:72:@30570.4]
  assign _T_60106 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11}; // @[Mux.scala 19:72:@30577.4]
  assign _T_60107 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,_T_60099}; // @[Mux.scala 19:72:@30578.4]
  assign _T_60109 = _T_2692 ? _T_60107 : 16'h0; // @[Mux.scala 19:72:@30579.4]
  assign _T_60116 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4}; // @[Mux.scala 19:72:@30586.4]
  assign _T_60123 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12}; // @[Mux.scala 19:72:@30593.4]
  assign _T_60124 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,_T_60116}; // @[Mux.scala 19:72:@30594.4]
  assign _T_60126 = _T_2693 ? _T_60124 : 16'h0; // @[Mux.scala 19:72:@30595.4]
  assign _T_60133 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5}; // @[Mux.scala 19:72:@30602.4]
  assign _T_60140 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13}; // @[Mux.scala 19:72:@30609.4]
  assign _T_60141 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,_T_60133}; // @[Mux.scala 19:72:@30610.4]
  assign _T_60143 = _T_2694 ? _T_60141 : 16'h0; // @[Mux.scala 19:72:@30611.4]
  assign _T_60150 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6}; // @[Mux.scala 19:72:@30618.4]
  assign _T_60157 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14}; // @[Mux.scala 19:72:@30625.4]
  assign _T_60158 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,_T_60150}; // @[Mux.scala 19:72:@30626.4]
  assign _T_60160 = _T_2695 ? _T_60158 : 16'h0; // @[Mux.scala 19:72:@30627.4]
  assign _T_60167 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7}; // @[Mux.scala 19:72:@30634.4]
  assign _T_60174 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15}; // @[Mux.scala 19:72:@30641.4]
  assign _T_60175 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,_T_60167}; // @[Mux.scala 19:72:@30642.4]
  assign _T_60177 = _T_2696 ? _T_60175 : 16'h0; // @[Mux.scala 19:72:@30643.4]
  assign _T_60192 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,_T_60055}; // @[Mux.scala 19:72:@30658.4]
  assign _T_60194 = _T_2697 ? _T_60192 : 16'h0; // @[Mux.scala 19:72:@30659.4]
  assign _T_60209 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,_T_60072}; // @[Mux.scala 19:72:@30674.4]
  assign _T_60211 = _T_2698 ? _T_60209 : 16'h0; // @[Mux.scala 19:72:@30675.4]
  assign _T_60226 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,_T_60089}; // @[Mux.scala 19:72:@30690.4]
  assign _T_60228 = _T_2699 ? _T_60226 : 16'h0; // @[Mux.scala 19:72:@30691.4]
  assign _T_60243 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,_T_60106}; // @[Mux.scala 19:72:@30706.4]
  assign _T_60245 = _T_2700 ? _T_60243 : 16'h0; // @[Mux.scala 19:72:@30707.4]
  assign _T_60260 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,_T_60123}; // @[Mux.scala 19:72:@30722.4]
  assign _T_60262 = _T_2701 ? _T_60260 : 16'h0; // @[Mux.scala 19:72:@30723.4]
  assign _T_60277 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,_T_60140}; // @[Mux.scala 19:72:@30738.4]
  assign _T_60279 = _T_2702 ? _T_60277 : 16'h0; // @[Mux.scala 19:72:@30739.4]
  assign _T_60294 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,_T_60157}; // @[Mux.scala 19:72:@30754.4]
  assign _T_60296 = _T_2703 ? _T_60294 : 16'h0; // @[Mux.scala 19:72:@30755.4]
  assign _T_60311 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,_T_60174}; // @[Mux.scala 19:72:@30770.4]
  assign _T_60313 = _T_2704 ? _T_60311 : 16'h0; // @[Mux.scala 19:72:@30771.4]
  assign _T_60314 = _T_60058 | _T_60075; // @[Mux.scala 19:72:@30772.4]
  assign _T_60315 = _T_60314 | _T_60092; // @[Mux.scala 19:72:@30773.4]
  assign _T_60316 = _T_60315 | _T_60109; // @[Mux.scala 19:72:@30774.4]
  assign _T_60317 = _T_60316 | _T_60126; // @[Mux.scala 19:72:@30775.4]
  assign _T_60318 = _T_60317 | _T_60143; // @[Mux.scala 19:72:@30776.4]
  assign _T_60319 = _T_60318 | _T_60160; // @[Mux.scala 19:72:@30777.4]
  assign _T_60320 = _T_60319 | _T_60177; // @[Mux.scala 19:72:@30778.4]
  assign _T_60321 = _T_60320 | _T_60194; // @[Mux.scala 19:72:@30779.4]
  assign _T_60322 = _T_60321 | _T_60211; // @[Mux.scala 19:72:@30780.4]
  assign _T_60323 = _T_60322 | _T_60228; // @[Mux.scala 19:72:@30781.4]
  assign _T_60324 = _T_60323 | _T_60245; // @[Mux.scala 19:72:@30782.4]
  assign _T_60325 = _T_60324 | _T_60262; // @[Mux.scala 19:72:@30783.4]
  assign _T_60326 = _T_60325 | _T_60279; // @[Mux.scala 19:72:@30784.4]
  assign _T_60327 = _T_60326 | _T_60296; // @[Mux.scala 19:72:@30785.4]
  assign _T_60328 = _T_60327 | _T_60313; // @[Mux.scala 19:72:@30786.4]
  assign _T_60906 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0}; // @[Mux.scala 19:72:@31136.4]
  assign _T_60913 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8}; // @[Mux.scala 19:72:@31143.4]
  assign _T_60914 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,_T_60906}; // @[Mux.scala 19:72:@31144.4]
  assign _T_60916 = _T_2689 ? _T_60914 : 16'h0; // @[Mux.scala 19:72:@31145.4]
  assign _T_60923 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1}; // @[Mux.scala 19:72:@31152.4]
  assign _T_60930 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9}; // @[Mux.scala 19:72:@31159.4]
  assign _T_60931 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,_T_60923}; // @[Mux.scala 19:72:@31160.4]
  assign _T_60933 = _T_2690 ? _T_60931 : 16'h0; // @[Mux.scala 19:72:@31161.4]
  assign _T_60940 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2}; // @[Mux.scala 19:72:@31168.4]
  assign _T_60947 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10}; // @[Mux.scala 19:72:@31175.4]
  assign _T_60948 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,_T_60940}; // @[Mux.scala 19:72:@31176.4]
  assign _T_60950 = _T_2691 ? _T_60948 : 16'h0; // @[Mux.scala 19:72:@31177.4]
  assign _T_60957 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3}; // @[Mux.scala 19:72:@31184.4]
  assign _T_60964 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11}; // @[Mux.scala 19:72:@31191.4]
  assign _T_60965 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,_T_60957}; // @[Mux.scala 19:72:@31192.4]
  assign _T_60967 = _T_2692 ? _T_60965 : 16'h0; // @[Mux.scala 19:72:@31193.4]
  assign _T_60974 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4}; // @[Mux.scala 19:72:@31200.4]
  assign _T_60981 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12}; // @[Mux.scala 19:72:@31207.4]
  assign _T_60982 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,_T_60974}; // @[Mux.scala 19:72:@31208.4]
  assign _T_60984 = _T_2693 ? _T_60982 : 16'h0; // @[Mux.scala 19:72:@31209.4]
  assign _T_60991 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5}; // @[Mux.scala 19:72:@31216.4]
  assign _T_60998 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13}; // @[Mux.scala 19:72:@31223.4]
  assign _T_60999 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,_T_60991}; // @[Mux.scala 19:72:@31224.4]
  assign _T_61001 = _T_2694 ? _T_60999 : 16'h0; // @[Mux.scala 19:72:@31225.4]
  assign _T_61008 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6}; // @[Mux.scala 19:72:@31232.4]
  assign _T_61015 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14}; // @[Mux.scala 19:72:@31239.4]
  assign _T_61016 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,_T_61008}; // @[Mux.scala 19:72:@31240.4]
  assign _T_61018 = _T_2695 ? _T_61016 : 16'h0; // @[Mux.scala 19:72:@31241.4]
  assign _T_61025 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7}; // @[Mux.scala 19:72:@31248.4]
  assign _T_61032 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15}; // @[Mux.scala 19:72:@31255.4]
  assign _T_61033 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,_T_61025}; // @[Mux.scala 19:72:@31256.4]
  assign _T_61035 = _T_2696 ? _T_61033 : 16'h0; // @[Mux.scala 19:72:@31257.4]
  assign _T_61050 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,_T_60913}; // @[Mux.scala 19:72:@31272.4]
  assign _T_61052 = _T_2697 ? _T_61050 : 16'h0; // @[Mux.scala 19:72:@31273.4]
  assign _T_61067 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,_T_60930}; // @[Mux.scala 19:72:@31288.4]
  assign _T_61069 = _T_2698 ? _T_61067 : 16'h0; // @[Mux.scala 19:72:@31289.4]
  assign _T_61084 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,_T_60947}; // @[Mux.scala 19:72:@31304.4]
  assign _T_61086 = _T_2699 ? _T_61084 : 16'h0; // @[Mux.scala 19:72:@31305.4]
  assign _T_61101 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,_T_60964}; // @[Mux.scala 19:72:@31320.4]
  assign _T_61103 = _T_2700 ? _T_61101 : 16'h0; // @[Mux.scala 19:72:@31321.4]
  assign _T_61118 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,_T_60981}; // @[Mux.scala 19:72:@31336.4]
  assign _T_61120 = _T_2701 ? _T_61118 : 16'h0; // @[Mux.scala 19:72:@31337.4]
  assign _T_61135 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,_T_60998}; // @[Mux.scala 19:72:@31352.4]
  assign _T_61137 = _T_2702 ? _T_61135 : 16'h0; // @[Mux.scala 19:72:@31353.4]
  assign _T_61152 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,_T_61015}; // @[Mux.scala 19:72:@31368.4]
  assign _T_61154 = _T_2703 ? _T_61152 : 16'h0; // @[Mux.scala 19:72:@31369.4]
  assign _T_61169 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,_T_61032}; // @[Mux.scala 19:72:@31384.4]
  assign _T_61171 = _T_2704 ? _T_61169 : 16'h0; // @[Mux.scala 19:72:@31385.4]
  assign _T_61172 = _T_60916 | _T_60933; // @[Mux.scala 19:72:@31386.4]
  assign _T_61173 = _T_61172 | _T_60950; // @[Mux.scala 19:72:@31387.4]
  assign _T_61174 = _T_61173 | _T_60967; // @[Mux.scala 19:72:@31388.4]
  assign _T_61175 = _T_61174 | _T_60984; // @[Mux.scala 19:72:@31389.4]
  assign _T_61176 = _T_61175 | _T_61001; // @[Mux.scala 19:72:@31390.4]
  assign _T_61177 = _T_61176 | _T_61018; // @[Mux.scala 19:72:@31391.4]
  assign _T_61178 = _T_61177 | _T_61035; // @[Mux.scala 19:72:@31392.4]
  assign _T_61179 = _T_61178 | _T_61052; // @[Mux.scala 19:72:@31393.4]
  assign _T_61180 = _T_61179 | _T_61069; // @[Mux.scala 19:72:@31394.4]
  assign _T_61181 = _T_61180 | _T_61086; // @[Mux.scala 19:72:@31395.4]
  assign _T_61182 = _T_61181 | _T_61103; // @[Mux.scala 19:72:@31396.4]
  assign _T_61183 = _T_61182 | _T_61120; // @[Mux.scala 19:72:@31397.4]
  assign _T_61184 = _T_61183 | _T_61137; // @[Mux.scala 19:72:@31398.4]
  assign _T_61185 = _T_61184 | _T_61154; // @[Mux.scala 19:72:@31399.4]
  assign _T_61186 = _T_61185 | _T_61171; // @[Mux.scala 19:72:@31400.4]
  assign _T_61764 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0}; // @[Mux.scala 19:72:@31750.4]
  assign _T_61771 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8}; // @[Mux.scala 19:72:@31757.4]
  assign _T_61772 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,_T_61764}; // @[Mux.scala 19:72:@31758.4]
  assign _T_61774 = _T_2689 ? _T_61772 : 16'h0; // @[Mux.scala 19:72:@31759.4]
  assign _T_61781 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1}; // @[Mux.scala 19:72:@31766.4]
  assign _T_61788 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9}; // @[Mux.scala 19:72:@31773.4]
  assign _T_61789 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,_T_61781}; // @[Mux.scala 19:72:@31774.4]
  assign _T_61791 = _T_2690 ? _T_61789 : 16'h0; // @[Mux.scala 19:72:@31775.4]
  assign _T_61798 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2}; // @[Mux.scala 19:72:@31782.4]
  assign _T_61805 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10}; // @[Mux.scala 19:72:@31789.4]
  assign _T_61806 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,_T_61798}; // @[Mux.scala 19:72:@31790.4]
  assign _T_61808 = _T_2691 ? _T_61806 : 16'h0; // @[Mux.scala 19:72:@31791.4]
  assign _T_61815 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3}; // @[Mux.scala 19:72:@31798.4]
  assign _T_61822 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11}; // @[Mux.scala 19:72:@31805.4]
  assign _T_61823 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,_T_61815}; // @[Mux.scala 19:72:@31806.4]
  assign _T_61825 = _T_2692 ? _T_61823 : 16'h0; // @[Mux.scala 19:72:@31807.4]
  assign _T_61832 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4}; // @[Mux.scala 19:72:@31814.4]
  assign _T_61839 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12}; // @[Mux.scala 19:72:@31821.4]
  assign _T_61840 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,_T_61832}; // @[Mux.scala 19:72:@31822.4]
  assign _T_61842 = _T_2693 ? _T_61840 : 16'h0; // @[Mux.scala 19:72:@31823.4]
  assign _T_61849 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5}; // @[Mux.scala 19:72:@31830.4]
  assign _T_61856 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13}; // @[Mux.scala 19:72:@31837.4]
  assign _T_61857 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,_T_61849}; // @[Mux.scala 19:72:@31838.4]
  assign _T_61859 = _T_2694 ? _T_61857 : 16'h0; // @[Mux.scala 19:72:@31839.4]
  assign _T_61866 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6}; // @[Mux.scala 19:72:@31846.4]
  assign _T_61873 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14}; // @[Mux.scala 19:72:@31853.4]
  assign _T_61874 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,_T_61866}; // @[Mux.scala 19:72:@31854.4]
  assign _T_61876 = _T_2695 ? _T_61874 : 16'h0; // @[Mux.scala 19:72:@31855.4]
  assign _T_61883 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7}; // @[Mux.scala 19:72:@31862.4]
  assign _T_61890 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15}; // @[Mux.scala 19:72:@31869.4]
  assign _T_61891 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,_T_61883}; // @[Mux.scala 19:72:@31870.4]
  assign _T_61893 = _T_2696 ? _T_61891 : 16'h0; // @[Mux.scala 19:72:@31871.4]
  assign _T_61908 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,_T_61771}; // @[Mux.scala 19:72:@31886.4]
  assign _T_61910 = _T_2697 ? _T_61908 : 16'h0; // @[Mux.scala 19:72:@31887.4]
  assign _T_61925 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,_T_61788}; // @[Mux.scala 19:72:@31902.4]
  assign _T_61927 = _T_2698 ? _T_61925 : 16'h0; // @[Mux.scala 19:72:@31903.4]
  assign _T_61942 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,_T_61805}; // @[Mux.scala 19:72:@31918.4]
  assign _T_61944 = _T_2699 ? _T_61942 : 16'h0; // @[Mux.scala 19:72:@31919.4]
  assign _T_61959 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,_T_61822}; // @[Mux.scala 19:72:@31934.4]
  assign _T_61961 = _T_2700 ? _T_61959 : 16'h0; // @[Mux.scala 19:72:@31935.4]
  assign _T_61976 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,_T_61839}; // @[Mux.scala 19:72:@31950.4]
  assign _T_61978 = _T_2701 ? _T_61976 : 16'h0; // @[Mux.scala 19:72:@31951.4]
  assign _T_61993 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,_T_61856}; // @[Mux.scala 19:72:@31966.4]
  assign _T_61995 = _T_2702 ? _T_61993 : 16'h0; // @[Mux.scala 19:72:@31967.4]
  assign _T_62010 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,_T_61873}; // @[Mux.scala 19:72:@31982.4]
  assign _T_62012 = _T_2703 ? _T_62010 : 16'h0; // @[Mux.scala 19:72:@31983.4]
  assign _T_62027 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,_T_61890}; // @[Mux.scala 19:72:@31998.4]
  assign _T_62029 = _T_2704 ? _T_62027 : 16'h0; // @[Mux.scala 19:72:@31999.4]
  assign _T_62030 = _T_61774 | _T_61791; // @[Mux.scala 19:72:@32000.4]
  assign _T_62031 = _T_62030 | _T_61808; // @[Mux.scala 19:72:@32001.4]
  assign _T_62032 = _T_62031 | _T_61825; // @[Mux.scala 19:72:@32002.4]
  assign _T_62033 = _T_62032 | _T_61842; // @[Mux.scala 19:72:@32003.4]
  assign _T_62034 = _T_62033 | _T_61859; // @[Mux.scala 19:72:@32004.4]
  assign _T_62035 = _T_62034 | _T_61876; // @[Mux.scala 19:72:@32005.4]
  assign _T_62036 = _T_62035 | _T_61893; // @[Mux.scala 19:72:@32006.4]
  assign _T_62037 = _T_62036 | _T_61910; // @[Mux.scala 19:72:@32007.4]
  assign _T_62038 = _T_62037 | _T_61927; // @[Mux.scala 19:72:@32008.4]
  assign _T_62039 = _T_62038 | _T_61944; // @[Mux.scala 19:72:@32009.4]
  assign _T_62040 = _T_62039 | _T_61961; // @[Mux.scala 19:72:@32010.4]
  assign _T_62041 = _T_62040 | _T_61978; // @[Mux.scala 19:72:@32011.4]
  assign _T_62042 = _T_62041 | _T_61995; // @[Mux.scala 19:72:@32012.4]
  assign _T_62043 = _T_62042 | _T_62012; // @[Mux.scala 19:72:@32013.4]
  assign _T_62044 = _T_62043 | _T_62029; // @[Mux.scala 19:72:@32014.4]
  assign _T_62622 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0}; // @[Mux.scala 19:72:@32364.4]
  assign _T_62629 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8}; // @[Mux.scala 19:72:@32371.4]
  assign _T_62630 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,_T_62622}; // @[Mux.scala 19:72:@32372.4]
  assign _T_62632 = _T_2689 ? _T_62630 : 16'h0; // @[Mux.scala 19:72:@32373.4]
  assign _T_62639 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1}; // @[Mux.scala 19:72:@32380.4]
  assign _T_62646 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9}; // @[Mux.scala 19:72:@32387.4]
  assign _T_62647 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,_T_62639}; // @[Mux.scala 19:72:@32388.4]
  assign _T_62649 = _T_2690 ? _T_62647 : 16'h0; // @[Mux.scala 19:72:@32389.4]
  assign _T_62656 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2}; // @[Mux.scala 19:72:@32396.4]
  assign _T_62663 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10}; // @[Mux.scala 19:72:@32403.4]
  assign _T_62664 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,_T_62656}; // @[Mux.scala 19:72:@32404.4]
  assign _T_62666 = _T_2691 ? _T_62664 : 16'h0; // @[Mux.scala 19:72:@32405.4]
  assign _T_62673 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3}; // @[Mux.scala 19:72:@32412.4]
  assign _T_62680 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11}; // @[Mux.scala 19:72:@32419.4]
  assign _T_62681 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,_T_62673}; // @[Mux.scala 19:72:@32420.4]
  assign _T_62683 = _T_2692 ? _T_62681 : 16'h0; // @[Mux.scala 19:72:@32421.4]
  assign _T_62690 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4}; // @[Mux.scala 19:72:@32428.4]
  assign _T_62697 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12}; // @[Mux.scala 19:72:@32435.4]
  assign _T_62698 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,_T_62690}; // @[Mux.scala 19:72:@32436.4]
  assign _T_62700 = _T_2693 ? _T_62698 : 16'h0; // @[Mux.scala 19:72:@32437.4]
  assign _T_62707 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5}; // @[Mux.scala 19:72:@32444.4]
  assign _T_62714 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13}; // @[Mux.scala 19:72:@32451.4]
  assign _T_62715 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,_T_62707}; // @[Mux.scala 19:72:@32452.4]
  assign _T_62717 = _T_2694 ? _T_62715 : 16'h0; // @[Mux.scala 19:72:@32453.4]
  assign _T_62724 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6}; // @[Mux.scala 19:72:@32460.4]
  assign _T_62731 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14}; // @[Mux.scala 19:72:@32467.4]
  assign _T_62732 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,_T_62724}; // @[Mux.scala 19:72:@32468.4]
  assign _T_62734 = _T_2695 ? _T_62732 : 16'h0; // @[Mux.scala 19:72:@32469.4]
  assign _T_62741 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7}; // @[Mux.scala 19:72:@32476.4]
  assign _T_62748 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15}; // @[Mux.scala 19:72:@32483.4]
  assign _T_62749 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,_T_62741}; // @[Mux.scala 19:72:@32484.4]
  assign _T_62751 = _T_2696 ? _T_62749 : 16'h0; // @[Mux.scala 19:72:@32485.4]
  assign _T_62766 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,_T_62629}; // @[Mux.scala 19:72:@32500.4]
  assign _T_62768 = _T_2697 ? _T_62766 : 16'h0; // @[Mux.scala 19:72:@32501.4]
  assign _T_62783 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,_T_62646}; // @[Mux.scala 19:72:@32516.4]
  assign _T_62785 = _T_2698 ? _T_62783 : 16'h0; // @[Mux.scala 19:72:@32517.4]
  assign _T_62800 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,_T_62663}; // @[Mux.scala 19:72:@32532.4]
  assign _T_62802 = _T_2699 ? _T_62800 : 16'h0; // @[Mux.scala 19:72:@32533.4]
  assign _T_62817 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,_T_62680}; // @[Mux.scala 19:72:@32548.4]
  assign _T_62819 = _T_2700 ? _T_62817 : 16'h0; // @[Mux.scala 19:72:@32549.4]
  assign _T_62834 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,_T_62697}; // @[Mux.scala 19:72:@32564.4]
  assign _T_62836 = _T_2701 ? _T_62834 : 16'h0; // @[Mux.scala 19:72:@32565.4]
  assign _T_62851 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,_T_62714}; // @[Mux.scala 19:72:@32580.4]
  assign _T_62853 = _T_2702 ? _T_62851 : 16'h0; // @[Mux.scala 19:72:@32581.4]
  assign _T_62868 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,_T_62731}; // @[Mux.scala 19:72:@32596.4]
  assign _T_62870 = _T_2703 ? _T_62868 : 16'h0; // @[Mux.scala 19:72:@32597.4]
  assign _T_62885 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,_T_62748}; // @[Mux.scala 19:72:@32612.4]
  assign _T_62887 = _T_2704 ? _T_62885 : 16'h0; // @[Mux.scala 19:72:@32613.4]
  assign _T_62888 = _T_62632 | _T_62649; // @[Mux.scala 19:72:@32614.4]
  assign _T_62889 = _T_62888 | _T_62666; // @[Mux.scala 19:72:@32615.4]
  assign _T_62890 = _T_62889 | _T_62683; // @[Mux.scala 19:72:@32616.4]
  assign _T_62891 = _T_62890 | _T_62700; // @[Mux.scala 19:72:@32617.4]
  assign _T_62892 = _T_62891 | _T_62717; // @[Mux.scala 19:72:@32618.4]
  assign _T_62893 = _T_62892 | _T_62734; // @[Mux.scala 19:72:@32619.4]
  assign _T_62894 = _T_62893 | _T_62751; // @[Mux.scala 19:72:@32620.4]
  assign _T_62895 = _T_62894 | _T_62768; // @[Mux.scala 19:72:@32621.4]
  assign _T_62896 = _T_62895 | _T_62785; // @[Mux.scala 19:72:@32622.4]
  assign _T_62897 = _T_62896 | _T_62802; // @[Mux.scala 19:72:@32623.4]
  assign _T_62898 = _T_62897 | _T_62819; // @[Mux.scala 19:72:@32624.4]
  assign _T_62899 = _T_62898 | _T_62836; // @[Mux.scala 19:72:@32625.4]
  assign _T_62900 = _T_62899 | _T_62853; // @[Mux.scala 19:72:@32626.4]
  assign _T_62901 = _T_62900 | _T_62870; // @[Mux.scala 19:72:@32627.4]
  assign _T_62902 = _T_62901 | _T_62887; // @[Mux.scala 19:72:@32628.4]
  assign _T_63480 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0}; // @[Mux.scala 19:72:@32978.4]
  assign _T_63487 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8}; // @[Mux.scala 19:72:@32985.4]
  assign _T_63488 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,_T_63480}; // @[Mux.scala 19:72:@32986.4]
  assign _T_63490 = _T_2689 ? _T_63488 : 16'h0; // @[Mux.scala 19:72:@32987.4]
  assign _T_63497 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1}; // @[Mux.scala 19:72:@32994.4]
  assign _T_63504 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9}; // @[Mux.scala 19:72:@33001.4]
  assign _T_63505 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,_T_63497}; // @[Mux.scala 19:72:@33002.4]
  assign _T_63507 = _T_2690 ? _T_63505 : 16'h0; // @[Mux.scala 19:72:@33003.4]
  assign _T_63514 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2}; // @[Mux.scala 19:72:@33010.4]
  assign _T_63521 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10}; // @[Mux.scala 19:72:@33017.4]
  assign _T_63522 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,_T_63514}; // @[Mux.scala 19:72:@33018.4]
  assign _T_63524 = _T_2691 ? _T_63522 : 16'h0; // @[Mux.scala 19:72:@33019.4]
  assign _T_63531 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3}; // @[Mux.scala 19:72:@33026.4]
  assign _T_63538 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11}; // @[Mux.scala 19:72:@33033.4]
  assign _T_63539 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,_T_63531}; // @[Mux.scala 19:72:@33034.4]
  assign _T_63541 = _T_2692 ? _T_63539 : 16'h0; // @[Mux.scala 19:72:@33035.4]
  assign _T_63548 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4}; // @[Mux.scala 19:72:@33042.4]
  assign _T_63555 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12}; // @[Mux.scala 19:72:@33049.4]
  assign _T_63556 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,_T_63548}; // @[Mux.scala 19:72:@33050.4]
  assign _T_63558 = _T_2693 ? _T_63556 : 16'h0; // @[Mux.scala 19:72:@33051.4]
  assign _T_63565 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5}; // @[Mux.scala 19:72:@33058.4]
  assign _T_63572 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13}; // @[Mux.scala 19:72:@33065.4]
  assign _T_63573 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,_T_63565}; // @[Mux.scala 19:72:@33066.4]
  assign _T_63575 = _T_2694 ? _T_63573 : 16'h0; // @[Mux.scala 19:72:@33067.4]
  assign _T_63582 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6}; // @[Mux.scala 19:72:@33074.4]
  assign _T_63589 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14}; // @[Mux.scala 19:72:@33081.4]
  assign _T_63590 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,_T_63582}; // @[Mux.scala 19:72:@33082.4]
  assign _T_63592 = _T_2695 ? _T_63590 : 16'h0; // @[Mux.scala 19:72:@33083.4]
  assign _T_63599 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7}; // @[Mux.scala 19:72:@33090.4]
  assign _T_63606 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15}; // @[Mux.scala 19:72:@33097.4]
  assign _T_63607 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,_T_63599}; // @[Mux.scala 19:72:@33098.4]
  assign _T_63609 = _T_2696 ? _T_63607 : 16'h0; // @[Mux.scala 19:72:@33099.4]
  assign _T_63624 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,_T_63487}; // @[Mux.scala 19:72:@33114.4]
  assign _T_63626 = _T_2697 ? _T_63624 : 16'h0; // @[Mux.scala 19:72:@33115.4]
  assign _T_63641 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,_T_63504}; // @[Mux.scala 19:72:@33130.4]
  assign _T_63643 = _T_2698 ? _T_63641 : 16'h0; // @[Mux.scala 19:72:@33131.4]
  assign _T_63658 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,_T_63521}; // @[Mux.scala 19:72:@33146.4]
  assign _T_63660 = _T_2699 ? _T_63658 : 16'h0; // @[Mux.scala 19:72:@33147.4]
  assign _T_63675 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,_T_63538}; // @[Mux.scala 19:72:@33162.4]
  assign _T_63677 = _T_2700 ? _T_63675 : 16'h0; // @[Mux.scala 19:72:@33163.4]
  assign _T_63692 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,_T_63555}; // @[Mux.scala 19:72:@33178.4]
  assign _T_63694 = _T_2701 ? _T_63692 : 16'h0; // @[Mux.scala 19:72:@33179.4]
  assign _T_63709 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,_T_63572}; // @[Mux.scala 19:72:@33194.4]
  assign _T_63711 = _T_2702 ? _T_63709 : 16'h0; // @[Mux.scala 19:72:@33195.4]
  assign _T_63726 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,_T_63589}; // @[Mux.scala 19:72:@33210.4]
  assign _T_63728 = _T_2703 ? _T_63726 : 16'h0; // @[Mux.scala 19:72:@33211.4]
  assign _T_63743 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,_T_63606}; // @[Mux.scala 19:72:@33226.4]
  assign _T_63745 = _T_2704 ? _T_63743 : 16'h0; // @[Mux.scala 19:72:@33227.4]
  assign _T_63746 = _T_63490 | _T_63507; // @[Mux.scala 19:72:@33228.4]
  assign _T_63747 = _T_63746 | _T_63524; // @[Mux.scala 19:72:@33229.4]
  assign _T_63748 = _T_63747 | _T_63541; // @[Mux.scala 19:72:@33230.4]
  assign _T_63749 = _T_63748 | _T_63558; // @[Mux.scala 19:72:@33231.4]
  assign _T_63750 = _T_63749 | _T_63575; // @[Mux.scala 19:72:@33232.4]
  assign _T_63751 = _T_63750 | _T_63592; // @[Mux.scala 19:72:@33233.4]
  assign _T_63752 = _T_63751 | _T_63609; // @[Mux.scala 19:72:@33234.4]
  assign _T_63753 = _T_63752 | _T_63626; // @[Mux.scala 19:72:@33235.4]
  assign _T_63754 = _T_63753 | _T_63643; // @[Mux.scala 19:72:@33236.4]
  assign _T_63755 = _T_63754 | _T_63660; // @[Mux.scala 19:72:@33237.4]
  assign _T_63756 = _T_63755 | _T_63677; // @[Mux.scala 19:72:@33238.4]
  assign _T_63757 = _T_63756 | _T_63694; // @[Mux.scala 19:72:@33239.4]
  assign _T_63758 = _T_63757 | _T_63711; // @[Mux.scala 19:72:@33240.4]
  assign _T_63759 = _T_63758 | _T_63728; // @[Mux.scala 19:72:@33241.4]
  assign _T_63760 = _T_63759 | _T_63745; // @[Mux.scala 19:72:@33242.4]
  assign _T_64338 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0}; // @[Mux.scala 19:72:@33592.4]
  assign _T_64345 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8}; // @[Mux.scala 19:72:@33599.4]
  assign _T_64346 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,_T_64338}; // @[Mux.scala 19:72:@33600.4]
  assign _T_64348 = _T_2689 ? _T_64346 : 16'h0; // @[Mux.scala 19:72:@33601.4]
  assign _T_64355 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1}; // @[Mux.scala 19:72:@33608.4]
  assign _T_64362 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9}; // @[Mux.scala 19:72:@33615.4]
  assign _T_64363 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,_T_64355}; // @[Mux.scala 19:72:@33616.4]
  assign _T_64365 = _T_2690 ? _T_64363 : 16'h0; // @[Mux.scala 19:72:@33617.4]
  assign _T_64372 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2}; // @[Mux.scala 19:72:@33624.4]
  assign _T_64379 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10}; // @[Mux.scala 19:72:@33631.4]
  assign _T_64380 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,_T_64372}; // @[Mux.scala 19:72:@33632.4]
  assign _T_64382 = _T_2691 ? _T_64380 : 16'h0; // @[Mux.scala 19:72:@33633.4]
  assign _T_64389 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3}; // @[Mux.scala 19:72:@33640.4]
  assign _T_64396 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11}; // @[Mux.scala 19:72:@33647.4]
  assign _T_64397 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,_T_64389}; // @[Mux.scala 19:72:@33648.4]
  assign _T_64399 = _T_2692 ? _T_64397 : 16'h0; // @[Mux.scala 19:72:@33649.4]
  assign _T_64406 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4}; // @[Mux.scala 19:72:@33656.4]
  assign _T_64413 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12}; // @[Mux.scala 19:72:@33663.4]
  assign _T_64414 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,_T_64406}; // @[Mux.scala 19:72:@33664.4]
  assign _T_64416 = _T_2693 ? _T_64414 : 16'h0; // @[Mux.scala 19:72:@33665.4]
  assign _T_64423 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5}; // @[Mux.scala 19:72:@33672.4]
  assign _T_64430 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13}; // @[Mux.scala 19:72:@33679.4]
  assign _T_64431 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,_T_64423}; // @[Mux.scala 19:72:@33680.4]
  assign _T_64433 = _T_2694 ? _T_64431 : 16'h0; // @[Mux.scala 19:72:@33681.4]
  assign _T_64440 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6}; // @[Mux.scala 19:72:@33688.4]
  assign _T_64447 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14}; // @[Mux.scala 19:72:@33695.4]
  assign _T_64448 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,_T_64440}; // @[Mux.scala 19:72:@33696.4]
  assign _T_64450 = _T_2695 ? _T_64448 : 16'h0; // @[Mux.scala 19:72:@33697.4]
  assign _T_64457 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7}; // @[Mux.scala 19:72:@33704.4]
  assign _T_64464 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15}; // @[Mux.scala 19:72:@33711.4]
  assign _T_64465 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,_T_64457}; // @[Mux.scala 19:72:@33712.4]
  assign _T_64467 = _T_2696 ? _T_64465 : 16'h0; // @[Mux.scala 19:72:@33713.4]
  assign _T_64482 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,_T_64345}; // @[Mux.scala 19:72:@33728.4]
  assign _T_64484 = _T_2697 ? _T_64482 : 16'h0; // @[Mux.scala 19:72:@33729.4]
  assign _T_64499 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,_T_64362}; // @[Mux.scala 19:72:@33744.4]
  assign _T_64501 = _T_2698 ? _T_64499 : 16'h0; // @[Mux.scala 19:72:@33745.4]
  assign _T_64516 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,_T_64379}; // @[Mux.scala 19:72:@33760.4]
  assign _T_64518 = _T_2699 ? _T_64516 : 16'h0; // @[Mux.scala 19:72:@33761.4]
  assign _T_64533 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,_T_64396}; // @[Mux.scala 19:72:@33776.4]
  assign _T_64535 = _T_2700 ? _T_64533 : 16'h0; // @[Mux.scala 19:72:@33777.4]
  assign _T_64550 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,_T_64413}; // @[Mux.scala 19:72:@33792.4]
  assign _T_64552 = _T_2701 ? _T_64550 : 16'h0; // @[Mux.scala 19:72:@33793.4]
  assign _T_64567 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,_T_64430}; // @[Mux.scala 19:72:@33808.4]
  assign _T_64569 = _T_2702 ? _T_64567 : 16'h0; // @[Mux.scala 19:72:@33809.4]
  assign _T_64584 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,_T_64447}; // @[Mux.scala 19:72:@33824.4]
  assign _T_64586 = _T_2703 ? _T_64584 : 16'h0; // @[Mux.scala 19:72:@33825.4]
  assign _T_64601 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,_T_64464}; // @[Mux.scala 19:72:@33840.4]
  assign _T_64603 = _T_2704 ? _T_64601 : 16'h0; // @[Mux.scala 19:72:@33841.4]
  assign _T_64604 = _T_64348 | _T_64365; // @[Mux.scala 19:72:@33842.4]
  assign _T_64605 = _T_64604 | _T_64382; // @[Mux.scala 19:72:@33843.4]
  assign _T_64606 = _T_64605 | _T_64399; // @[Mux.scala 19:72:@33844.4]
  assign _T_64607 = _T_64606 | _T_64416; // @[Mux.scala 19:72:@33845.4]
  assign _T_64608 = _T_64607 | _T_64433; // @[Mux.scala 19:72:@33846.4]
  assign _T_64609 = _T_64608 | _T_64450; // @[Mux.scala 19:72:@33847.4]
  assign _T_64610 = _T_64609 | _T_64467; // @[Mux.scala 19:72:@33848.4]
  assign _T_64611 = _T_64610 | _T_64484; // @[Mux.scala 19:72:@33849.4]
  assign _T_64612 = _T_64611 | _T_64501; // @[Mux.scala 19:72:@33850.4]
  assign _T_64613 = _T_64612 | _T_64518; // @[Mux.scala 19:72:@33851.4]
  assign _T_64614 = _T_64613 | _T_64535; // @[Mux.scala 19:72:@33852.4]
  assign _T_64615 = _T_64614 | _T_64552; // @[Mux.scala 19:72:@33853.4]
  assign _T_64616 = _T_64615 | _T_64569; // @[Mux.scala 19:72:@33854.4]
  assign _T_64617 = _T_64616 | _T_64586; // @[Mux.scala 19:72:@33855.4]
  assign _T_64618 = _T_64617 | _T_64603; // @[Mux.scala 19:72:@33856.4]
  assign _T_65196 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0}; // @[Mux.scala 19:72:@34206.4]
  assign _T_65203 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8}; // @[Mux.scala 19:72:@34213.4]
  assign _T_65204 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,_T_65196}; // @[Mux.scala 19:72:@34214.4]
  assign _T_65206 = _T_2689 ? _T_65204 : 16'h0; // @[Mux.scala 19:72:@34215.4]
  assign _T_65213 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1}; // @[Mux.scala 19:72:@34222.4]
  assign _T_65220 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9}; // @[Mux.scala 19:72:@34229.4]
  assign _T_65221 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,_T_65213}; // @[Mux.scala 19:72:@34230.4]
  assign _T_65223 = _T_2690 ? _T_65221 : 16'h0; // @[Mux.scala 19:72:@34231.4]
  assign _T_65230 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2}; // @[Mux.scala 19:72:@34238.4]
  assign _T_65237 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10}; // @[Mux.scala 19:72:@34245.4]
  assign _T_65238 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,_T_65230}; // @[Mux.scala 19:72:@34246.4]
  assign _T_65240 = _T_2691 ? _T_65238 : 16'h0; // @[Mux.scala 19:72:@34247.4]
  assign _T_65247 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3}; // @[Mux.scala 19:72:@34254.4]
  assign _T_65254 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11}; // @[Mux.scala 19:72:@34261.4]
  assign _T_65255 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,_T_65247}; // @[Mux.scala 19:72:@34262.4]
  assign _T_65257 = _T_2692 ? _T_65255 : 16'h0; // @[Mux.scala 19:72:@34263.4]
  assign _T_65264 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4}; // @[Mux.scala 19:72:@34270.4]
  assign _T_65271 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12}; // @[Mux.scala 19:72:@34277.4]
  assign _T_65272 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,_T_65264}; // @[Mux.scala 19:72:@34278.4]
  assign _T_65274 = _T_2693 ? _T_65272 : 16'h0; // @[Mux.scala 19:72:@34279.4]
  assign _T_65281 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5}; // @[Mux.scala 19:72:@34286.4]
  assign _T_65288 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13}; // @[Mux.scala 19:72:@34293.4]
  assign _T_65289 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,_T_65281}; // @[Mux.scala 19:72:@34294.4]
  assign _T_65291 = _T_2694 ? _T_65289 : 16'h0; // @[Mux.scala 19:72:@34295.4]
  assign _T_65298 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6}; // @[Mux.scala 19:72:@34302.4]
  assign _T_65305 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14}; // @[Mux.scala 19:72:@34309.4]
  assign _T_65306 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,_T_65298}; // @[Mux.scala 19:72:@34310.4]
  assign _T_65308 = _T_2695 ? _T_65306 : 16'h0; // @[Mux.scala 19:72:@34311.4]
  assign _T_65315 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7}; // @[Mux.scala 19:72:@34318.4]
  assign _T_65322 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15}; // @[Mux.scala 19:72:@34325.4]
  assign _T_65323 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,_T_65315}; // @[Mux.scala 19:72:@34326.4]
  assign _T_65325 = _T_2696 ? _T_65323 : 16'h0; // @[Mux.scala 19:72:@34327.4]
  assign _T_65340 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,_T_65203}; // @[Mux.scala 19:72:@34342.4]
  assign _T_65342 = _T_2697 ? _T_65340 : 16'h0; // @[Mux.scala 19:72:@34343.4]
  assign _T_65357 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,_T_65220}; // @[Mux.scala 19:72:@34358.4]
  assign _T_65359 = _T_2698 ? _T_65357 : 16'h0; // @[Mux.scala 19:72:@34359.4]
  assign _T_65374 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,_T_65237}; // @[Mux.scala 19:72:@34374.4]
  assign _T_65376 = _T_2699 ? _T_65374 : 16'h0; // @[Mux.scala 19:72:@34375.4]
  assign _T_65391 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,_T_65254}; // @[Mux.scala 19:72:@34390.4]
  assign _T_65393 = _T_2700 ? _T_65391 : 16'h0; // @[Mux.scala 19:72:@34391.4]
  assign _T_65408 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,_T_65271}; // @[Mux.scala 19:72:@34406.4]
  assign _T_65410 = _T_2701 ? _T_65408 : 16'h0; // @[Mux.scala 19:72:@34407.4]
  assign _T_65425 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,_T_65288}; // @[Mux.scala 19:72:@34422.4]
  assign _T_65427 = _T_2702 ? _T_65425 : 16'h0; // @[Mux.scala 19:72:@34423.4]
  assign _T_65442 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,_T_65305}; // @[Mux.scala 19:72:@34438.4]
  assign _T_65444 = _T_2703 ? _T_65442 : 16'h0; // @[Mux.scala 19:72:@34439.4]
  assign _T_65459 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,_T_65322}; // @[Mux.scala 19:72:@34454.4]
  assign _T_65461 = _T_2704 ? _T_65459 : 16'h0; // @[Mux.scala 19:72:@34455.4]
  assign _T_65462 = _T_65206 | _T_65223; // @[Mux.scala 19:72:@34456.4]
  assign _T_65463 = _T_65462 | _T_65240; // @[Mux.scala 19:72:@34457.4]
  assign _T_65464 = _T_65463 | _T_65257; // @[Mux.scala 19:72:@34458.4]
  assign _T_65465 = _T_65464 | _T_65274; // @[Mux.scala 19:72:@34459.4]
  assign _T_65466 = _T_65465 | _T_65291; // @[Mux.scala 19:72:@34460.4]
  assign _T_65467 = _T_65466 | _T_65308; // @[Mux.scala 19:72:@34461.4]
  assign _T_65468 = _T_65467 | _T_65325; // @[Mux.scala 19:72:@34462.4]
  assign _T_65469 = _T_65468 | _T_65342; // @[Mux.scala 19:72:@34463.4]
  assign _T_65470 = _T_65469 | _T_65359; // @[Mux.scala 19:72:@34464.4]
  assign _T_65471 = _T_65470 | _T_65376; // @[Mux.scala 19:72:@34465.4]
  assign _T_65472 = _T_65471 | _T_65393; // @[Mux.scala 19:72:@34466.4]
  assign _T_65473 = _T_65472 | _T_65410; // @[Mux.scala 19:72:@34467.4]
  assign _T_65474 = _T_65473 | _T_65427; // @[Mux.scala 19:72:@34468.4]
  assign _T_65475 = _T_65474 | _T_65444; // @[Mux.scala 19:72:@34469.4]
  assign _T_65476 = _T_65475 | _T_65461; // @[Mux.scala 19:72:@34470.4]
  assign _T_88268 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[LoadQueue.scala 191:60:@35143.4]
  assign _T_88269 = conflictPReg_0_3 ? 2'h3 : _T_88268; // @[LoadQueue.scala 191:60:@35144.4]
  assign _T_88270 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_88269}; // @[LoadQueue.scala 191:60:@35145.4]
  assign _T_88271 = conflictPReg_0_5 ? 3'h5 : _T_88270; // @[LoadQueue.scala 191:60:@35146.4]
  assign _T_88272 = conflictPReg_0_6 ? 3'h6 : _T_88271; // @[LoadQueue.scala 191:60:@35147.4]
  assign _T_88273 = conflictPReg_0_7 ? 3'h7 : _T_88272; // @[LoadQueue.scala 191:60:@35148.4]
  assign _T_88274 = conflictPReg_0_8 ? 4'h8 : {{1'd0}, _T_88273}; // @[LoadQueue.scala 191:60:@35149.4]
  assign _T_88275 = conflictPReg_0_9 ? 4'h9 : _T_88274; // @[LoadQueue.scala 191:60:@35150.4]
  assign _T_88276 = conflictPReg_0_10 ? 4'ha : _T_88275; // @[LoadQueue.scala 191:60:@35151.4]
  assign _T_88277 = conflictPReg_0_11 ? 4'hb : _T_88276; // @[LoadQueue.scala 191:60:@35152.4]
  assign _T_88278 = conflictPReg_0_12 ? 4'hc : _T_88277; // @[LoadQueue.scala 191:60:@35153.4]
  assign _T_88279 = conflictPReg_0_13 ? 4'hd : _T_88278; // @[LoadQueue.scala 191:60:@35154.4]
  assign _T_88280 = conflictPReg_0_14 ? 4'he : _T_88279; // @[LoadQueue.scala 191:60:@35155.4]
  assign _T_88281 = conflictPReg_0_15 ? 4'hf : _T_88280; // @[LoadQueue.scala 191:60:@35156.4]
  assign _T_88284 = conflictPReg_0_0 | conflictPReg_0_1; // @[LoadQueue.scala 192:43:@35158.4]
  assign _T_88285 = _T_88284 | conflictPReg_0_2; // @[LoadQueue.scala 192:43:@35159.4]
  assign _T_88286 = _T_88285 | conflictPReg_0_3; // @[LoadQueue.scala 192:43:@35160.4]
  assign _T_88287 = _T_88286 | conflictPReg_0_4; // @[LoadQueue.scala 192:43:@35161.4]
  assign _T_88288 = _T_88287 | conflictPReg_0_5; // @[LoadQueue.scala 192:43:@35162.4]
  assign _T_88289 = _T_88288 | conflictPReg_0_6; // @[LoadQueue.scala 192:43:@35163.4]
  assign _T_88290 = _T_88289 | conflictPReg_0_7; // @[LoadQueue.scala 192:43:@35164.4]
  assign _T_88291 = _T_88290 | conflictPReg_0_8; // @[LoadQueue.scala 192:43:@35165.4]
  assign _T_88292 = _T_88291 | conflictPReg_0_9; // @[LoadQueue.scala 192:43:@35166.4]
  assign _T_88293 = _T_88292 | conflictPReg_0_10; // @[LoadQueue.scala 192:43:@35167.4]
  assign _T_88294 = _T_88293 | conflictPReg_0_11; // @[LoadQueue.scala 192:43:@35168.4]
  assign _T_88295 = _T_88294 | conflictPReg_0_12; // @[LoadQueue.scala 192:43:@35169.4]
  assign _T_88296 = _T_88295 | conflictPReg_0_13; // @[LoadQueue.scala 192:43:@35170.4]
  assign _T_88297 = _T_88296 | conflictPReg_0_14; // @[LoadQueue.scala 192:43:@35171.4]
  assign _T_88298 = _T_88297 | conflictPReg_0_15; // @[LoadQueue.scala 192:43:@35172.4]
  assign _GEN_864 = 4'h0 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_865 = 4'h1 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_866 = 4'h2 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_867 = 4'h3 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_868 = 4'h4 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_869 = 4'h5 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_870 = 4'h6 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_871 = 4'h7 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_872 = 4'h8 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_873 = 4'h9 == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_874 = 4'ha == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_875 = 4'hb == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_876 = 4'hc == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_877 = 4'hd == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_878 = 4'he == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_879 = 4'hf == _T_88281; // @[LoadQueue.scala 193:43:@35174.6]
  assign _GEN_881 = 4'h1 == _T_88281 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_882 = 4'h2 == _T_88281 ? shiftedStoreDataKnownPReg_2 : _GEN_881; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_883 = 4'h3 == _T_88281 ? shiftedStoreDataKnownPReg_3 : _GEN_882; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_884 = 4'h4 == _T_88281 ? shiftedStoreDataKnownPReg_4 : _GEN_883; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_885 = 4'h5 == _T_88281 ? shiftedStoreDataKnownPReg_5 : _GEN_884; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_886 = 4'h6 == _T_88281 ? shiftedStoreDataKnownPReg_6 : _GEN_885; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_887 = 4'h7 == _T_88281 ? shiftedStoreDataKnownPReg_7 : _GEN_886; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_888 = 4'h8 == _T_88281 ? shiftedStoreDataKnownPReg_8 : _GEN_887; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_889 = 4'h9 == _T_88281 ? shiftedStoreDataKnownPReg_9 : _GEN_888; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_890 = 4'ha == _T_88281 ? shiftedStoreDataKnownPReg_10 : _GEN_889; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_891 = 4'hb == _T_88281 ? shiftedStoreDataKnownPReg_11 : _GEN_890; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_892 = 4'hc == _T_88281 ? shiftedStoreDataKnownPReg_12 : _GEN_891; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_893 = 4'hd == _T_88281 ? shiftedStoreDataKnownPReg_13 : _GEN_892; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_894 = 4'he == _T_88281 ? shiftedStoreDataKnownPReg_14 : _GEN_893; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_895 = 4'hf == _T_88281 ? shiftedStoreDataKnownPReg_15 : _GEN_894; // @[LoadQueue.scala 194:31:@35175.6]
  assign _GEN_897 = 4'h1 == _T_88281 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_898 = 4'h2 == _T_88281 ? shiftedStoreDataQPreg_2 : _GEN_897; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_899 = 4'h3 == _T_88281 ? shiftedStoreDataQPreg_3 : _GEN_898; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_900 = 4'h4 == _T_88281 ? shiftedStoreDataQPreg_4 : _GEN_899; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_901 = 4'h5 == _T_88281 ? shiftedStoreDataQPreg_5 : _GEN_900; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_902 = 4'h6 == _T_88281 ? shiftedStoreDataQPreg_6 : _GEN_901; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_903 = 4'h7 == _T_88281 ? shiftedStoreDataQPreg_7 : _GEN_902; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_904 = 4'h8 == _T_88281 ? shiftedStoreDataQPreg_8 : _GEN_903; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_905 = 4'h9 == _T_88281 ? shiftedStoreDataQPreg_9 : _GEN_904; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_906 = 4'ha == _T_88281 ? shiftedStoreDataQPreg_10 : _GEN_905; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_907 = 4'hb == _T_88281 ? shiftedStoreDataQPreg_11 : _GEN_906; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_908 = 4'hc == _T_88281 ? shiftedStoreDataQPreg_12 : _GEN_907; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_909 = 4'hd == _T_88281 ? shiftedStoreDataQPreg_13 : _GEN_908; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_910 = 4'he == _T_88281 ? shiftedStoreDataQPreg_14 : _GEN_909; // @[LoadQueue.scala 195:31:@35176.6]
  assign _GEN_911 = 4'hf == _T_88281 ? shiftedStoreDataQPreg_15 : _GEN_910; // @[LoadQueue.scala 195:31:@35176.6]
  assign lastConflict_0_0 = _T_88298 ? _GEN_864 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_1 = _T_88298 ? _GEN_865 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_2 = _T_88298 ? _GEN_866 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_3 = _T_88298 ? _GEN_867 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_4 = _T_88298 ? _GEN_868 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_5 = _T_88298 ? _GEN_869 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_6 = _T_88298 ? _GEN_870 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_7 = _T_88298 ? _GEN_871 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_8 = _T_88298 ? _GEN_872 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_9 = _T_88298 ? _GEN_873 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_10 = _T_88298 ? _GEN_874 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_11 = _T_88298 ? _GEN_875 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_12 = _T_88298 ? _GEN_876 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_13 = _T_88298 ? _GEN_877 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_14 = _T_88298 ? _GEN_878 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign lastConflict_0_15 = _T_88298 ? _GEN_879 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign canBypass_0 = _T_88298 ? _GEN_895 : 1'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign bypassVal_0 = _T_88298 ? _GEN_911 : 32'h0; // @[LoadQueue.scala 192:53:@35173.4]
  assign _T_88404 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[LoadQueue.scala 191:60:@35230.4]
  assign _T_88405 = conflictPReg_1_3 ? 2'h3 : _T_88404; // @[LoadQueue.scala 191:60:@35231.4]
  assign _T_88406 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_88405}; // @[LoadQueue.scala 191:60:@35232.4]
  assign _T_88407 = conflictPReg_1_5 ? 3'h5 : _T_88406; // @[LoadQueue.scala 191:60:@35233.4]
  assign _T_88408 = conflictPReg_1_6 ? 3'h6 : _T_88407; // @[LoadQueue.scala 191:60:@35234.4]
  assign _T_88409 = conflictPReg_1_7 ? 3'h7 : _T_88408; // @[LoadQueue.scala 191:60:@35235.4]
  assign _T_88410 = conflictPReg_1_8 ? 4'h8 : {{1'd0}, _T_88409}; // @[LoadQueue.scala 191:60:@35236.4]
  assign _T_88411 = conflictPReg_1_9 ? 4'h9 : _T_88410; // @[LoadQueue.scala 191:60:@35237.4]
  assign _T_88412 = conflictPReg_1_10 ? 4'ha : _T_88411; // @[LoadQueue.scala 191:60:@35238.4]
  assign _T_88413 = conflictPReg_1_11 ? 4'hb : _T_88412; // @[LoadQueue.scala 191:60:@35239.4]
  assign _T_88414 = conflictPReg_1_12 ? 4'hc : _T_88413; // @[LoadQueue.scala 191:60:@35240.4]
  assign _T_88415 = conflictPReg_1_13 ? 4'hd : _T_88414; // @[LoadQueue.scala 191:60:@35241.4]
  assign _T_88416 = conflictPReg_1_14 ? 4'he : _T_88415; // @[LoadQueue.scala 191:60:@35242.4]
  assign _T_88417 = conflictPReg_1_15 ? 4'hf : _T_88416; // @[LoadQueue.scala 191:60:@35243.4]
  assign _T_88420 = conflictPReg_1_0 | conflictPReg_1_1; // @[LoadQueue.scala 192:43:@35245.4]
  assign _T_88421 = _T_88420 | conflictPReg_1_2; // @[LoadQueue.scala 192:43:@35246.4]
  assign _T_88422 = _T_88421 | conflictPReg_1_3; // @[LoadQueue.scala 192:43:@35247.4]
  assign _T_88423 = _T_88422 | conflictPReg_1_4; // @[LoadQueue.scala 192:43:@35248.4]
  assign _T_88424 = _T_88423 | conflictPReg_1_5; // @[LoadQueue.scala 192:43:@35249.4]
  assign _T_88425 = _T_88424 | conflictPReg_1_6; // @[LoadQueue.scala 192:43:@35250.4]
  assign _T_88426 = _T_88425 | conflictPReg_1_7; // @[LoadQueue.scala 192:43:@35251.4]
  assign _T_88427 = _T_88426 | conflictPReg_1_8; // @[LoadQueue.scala 192:43:@35252.4]
  assign _T_88428 = _T_88427 | conflictPReg_1_9; // @[LoadQueue.scala 192:43:@35253.4]
  assign _T_88429 = _T_88428 | conflictPReg_1_10; // @[LoadQueue.scala 192:43:@35254.4]
  assign _T_88430 = _T_88429 | conflictPReg_1_11; // @[LoadQueue.scala 192:43:@35255.4]
  assign _T_88431 = _T_88430 | conflictPReg_1_12; // @[LoadQueue.scala 192:43:@35256.4]
  assign _T_88432 = _T_88431 | conflictPReg_1_13; // @[LoadQueue.scala 192:43:@35257.4]
  assign _T_88433 = _T_88432 | conflictPReg_1_14; // @[LoadQueue.scala 192:43:@35258.4]
  assign _T_88434 = _T_88433 | conflictPReg_1_15; // @[LoadQueue.scala 192:43:@35259.4]
  assign _GEN_930 = 4'h0 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_931 = 4'h1 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_932 = 4'h2 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_933 = 4'h3 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_934 = 4'h4 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_935 = 4'h5 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_936 = 4'h6 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_937 = 4'h7 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_938 = 4'h8 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_939 = 4'h9 == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_940 = 4'ha == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_941 = 4'hb == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_942 = 4'hc == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_943 = 4'hd == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_944 = 4'he == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_945 = 4'hf == _T_88417; // @[LoadQueue.scala 193:43:@35261.6]
  assign _GEN_947 = 4'h1 == _T_88417 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_948 = 4'h2 == _T_88417 ? shiftedStoreDataKnownPReg_2 : _GEN_947; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_949 = 4'h3 == _T_88417 ? shiftedStoreDataKnownPReg_3 : _GEN_948; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_950 = 4'h4 == _T_88417 ? shiftedStoreDataKnownPReg_4 : _GEN_949; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_951 = 4'h5 == _T_88417 ? shiftedStoreDataKnownPReg_5 : _GEN_950; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_952 = 4'h6 == _T_88417 ? shiftedStoreDataKnownPReg_6 : _GEN_951; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_953 = 4'h7 == _T_88417 ? shiftedStoreDataKnownPReg_7 : _GEN_952; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_954 = 4'h8 == _T_88417 ? shiftedStoreDataKnownPReg_8 : _GEN_953; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_955 = 4'h9 == _T_88417 ? shiftedStoreDataKnownPReg_9 : _GEN_954; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_956 = 4'ha == _T_88417 ? shiftedStoreDataKnownPReg_10 : _GEN_955; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_957 = 4'hb == _T_88417 ? shiftedStoreDataKnownPReg_11 : _GEN_956; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_958 = 4'hc == _T_88417 ? shiftedStoreDataKnownPReg_12 : _GEN_957; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_959 = 4'hd == _T_88417 ? shiftedStoreDataKnownPReg_13 : _GEN_958; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_960 = 4'he == _T_88417 ? shiftedStoreDataKnownPReg_14 : _GEN_959; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_961 = 4'hf == _T_88417 ? shiftedStoreDataKnownPReg_15 : _GEN_960; // @[LoadQueue.scala 194:31:@35262.6]
  assign _GEN_963 = 4'h1 == _T_88417 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_964 = 4'h2 == _T_88417 ? shiftedStoreDataQPreg_2 : _GEN_963; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_965 = 4'h3 == _T_88417 ? shiftedStoreDataQPreg_3 : _GEN_964; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_966 = 4'h4 == _T_88417 ? shiftedStoreDataQPreg_4 : _GEN_965; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_967 = 4'h5 == _T_88417 ? shiftedStoreDataQPreg_5 : _GEN_966; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_968 = 4'h6 == _T_88417 ? shiftedStoreDataQPreg_6 : _GEN_967; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_969 = 4'h7 == _T_88417 ? shiftedStoreDataQPreg_7 : _GEN_968; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_970 = 4'h8 == _T_88417 ? shiftedStoreDataQPreg_8 : _GEN_969; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_971 = 4'h9 == _T_88417 ? shiftedStoreDataQPreg_9 : _GEN_970; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_972 = 4'ha == _T_88417 ? shiftedStoreDataQPreg_10 : _GEN_971; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_973 = 4'hb == _T_88417 ? shiftedStoreDataQPreg_11 : _GEN_972; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_974 = 4'hc == _T_88417 ? shiftedStoreDataQPreg_12 : _GEN_973; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_975 = 4'hd == _T_88417 ? shiftedStoreDataQPreg_13 : _GEN_974; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_976 = 4'he == _T_88417 ? shiftedStoreDataQPreg_14 : _GEN_975; // @[LoadQueue.scala 195:31:@35263.6]
  assign _GEN_977 = 4'hf == _T_88417 ? shiftedStoreDataQPreg_15 : _GEN_976; // @[LoadQueue.scala 195:31:@35263.6]
  assign lastConflict_1_0 = _T_88434 ? _GEN_930 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_1 = _T_88434 ? _GEN_931 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_2 = _T_88434 ? _GEN_932 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_3 = _T_88434 ? _GEN_933 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_4 = _T_88434 ? _GEN_934 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_5 = _T_88434 ? _GEN_935 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_6 = _T_88434 ? _GEN_936 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_7 = _T_88434 ? _GEN_937 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_8 = _T_88434 ? _GEN_938 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_9 = _T_88434 ? _GEN_939 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_10 = _T_88434 ? _GEN_940 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_11 = _T_88434 ? _GEN_941 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_12 = _T_88434 ? _GEN_942 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_13 = _T_88434 ? _GEN_943 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_14 = _T_88434 ? _GEN_944 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign lastConflict_1_15 = _T_88434 ? _GEN_945 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign canBypass_1 = _T_88434 ? _GEN_961 : 1'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign bypassVal_1 = _T_88434 ? _GEN_977 : 32'h0; // @[LoadQueue.scala 192:53:@35260.4]
  assign _T_88540 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[LoadQueue.scala 191:60:@35317.4]
  assign _T_88541 = conflictPReg_2_3 ? 2'h3 : _T_88540; // @[LoadQueue.scala 191:60:@35318.4]
  assign _T_88542 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_88541}; // @[LoadQueue.scala 191:60:@35319.4]
  assign _T_88543 = conflictPReg_2_5 ? 3'h5 : _T_88542; // @[LoadQueue.scala 191:60:@35320.4]
  assign _T_88544 = conflictPReg_2_6 ? 3'h6 : _T_88543; // @[LoadQueue.scala 191:60:@35321.4]
  assign _T_88545 = conflictPReg_2_7 ? 3'h7 : _T_88544; // @[LoadQueue.scala 191:60:@35322.4]
  assign _T_88546 = conflictPReg_2_8 ? 4'h8 : {{1'd0}, _T_88545}; // @[LoadQueue.scala 191:60:@35323.4]
  assign _T_88547 = conflictPReg_2_9 ? 4'h9 : _T_88546; // @[LoadQueue.scala 191:60:@35324.4]
  assign _T_88548 = conflictPReg_2_10 ? 4'ha : _T_88547; // @[LoadQueue.scala 191:60:@35325.4]
  assign _T_88549 = conflictPReg_2_11 ? 4'hb : _T_88548; // @[LoadQueue.scala 191:60:@35326.4]
  assign _T_88550 = conflictPReg_2_12 ? 4'hc : _T_88549; // @[LoadQueue.scala 191:60:@35327.4]
  assign _T_88551 = conflictPReg_2_13 ? 4'hd : _T_88550; // @[LoadQueue.scala 191:60:@35328.4]
  assign _T_88552 = conflictPReg_2_14 ? 4'he : _T_88551; // @[LoadQueue.scala 191:60:@35329.4]
  assign _T_88553 = conflictPReg_2_15 ? 4'hf : _T_88552; // @[LoadQueue.scala 191:60:@35330.4]
  assign _T_88556 = conflictPReg_2_0 | conflictPReg_2_1; // @[LoadQueue.scala 192:43:@35332.4]
  assign _T_88557 = _T_88556 | conflictPReg_2_2; // @[LoadQueue.scala 192:43:@35333.4]
  assign _T_88558 = _T_88557 | conflictPReg_2_3; // @[LoadQueue.scala 192:43:@35334.4]
  assign _T_88559 = _T_88558 | conflictPReg_2_4; // @[LoadQueue.scala 192:43:@35335.4]
  assign _T_88560 = _T_88559 | conflictPReg_2_5; // @[LoadQueue.scala 192:43:@35336.4]
  assign _T_88561 = _T_88560 | conflictPReg_2_6; // @[LoadQueue.scala 192:43:@35337.4]
  assign _T_88562 = _T_88561 | conflictPReg_2_7; // @[LoadQueue.scala 192:43:@35338.4]
  assign _T_88563 = _T_88562 | conflictPReg_2_8; // @[LoadQueue.scala 192:43:@35339.4]
  assign _T_88564 = _T_88563 | conflictPReg_2_9; // @[LoadQueue.scala 192:43:@35340.4]
  assign _T_88565 = _T_88564 | conflictPReg_2_10; // @[LoadQueue.scala 192:43:@35341.4]
  assign _T_88566 = _T_88565 | conflictPReg_2_11; // @[LoadQueue.scala 192:43:@35342.4]
  assign _T_88567 = _T_88566 | conflictPReg_2_12; // @[LoadQueue.scala 192:43:@35343.4]
  assign _T_88568 = _T_88567 | conflictPReg_2_13; // @[LoadQueue.scala 192:43:@35344.4]
  assign _T_88569 = _T_88568 | conflictPReg_2_14; // @[LoadQueue.scala 192:43:@35345.4]
  assign _T_88570 = _T_88569 | conflictPReg_2_15; // @[LoadQueue.scala 192:43:@35346.4]
  assign _GEN_996 = 4'h0 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_997 = 4'h1 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_998 = 4'h2 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_999 = 4'h3 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1000 = 4'h4 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1001 = 4'h5 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1002 = 4'h6 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1003 = 4'h7 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1004 = 4'h8 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1005 = 4'h9 == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1006 = 4'ha == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1007 = 4'hb == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1008 = 4'hc == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1009 = 4'hd == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1010 = 4'he == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1011 = 4'hf == _T_88553; // @[LoadQueue.scala 193:43:@35348.6]
  assign _GEN_1013 = 4'h1 == _T_88553 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1014 = 4'h2 == _T_88553 ? shiftedStoreDataKnownPReg_2 : _GEN_1013; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1015 = 4'h3 == _T_88553 ? shiftedStoreDataKnownPReg_3 : _GEN_1014; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1016 = 4'h4 == _T_88553 ? shiftedStoreDataKnownPReg_4 : _GEN_1015; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1017 = 4'h5 == _T_88553 ? shiftedStoreDataKnownPReg_5 : _GEN_1016; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1018 = 4'h6 == _T_88553 ? shiftedStoreDataKnownPReg_6 : _GEN_1017; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1019 = 4'h7 == _T_88553 ? shiftedStoreDataKnownPReg_7 : _GEN_1018; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1020 = 4'h8 == _T_88553 ? shiftedStoreDataKnownPReg_8 : _GEN_1019; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1021 = 4'h9 == _T_88553 ? shiftedStoreDataKnownPReg_9 : _GEN_1020; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1022 = 4'ha == _T_88553 ? shiftedStoreDataKnownPReg_10 : _GEN_1021; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1023 = 4'hb == _T_88553 ? shiftedStoreDataKnownPReg_11 : _GEN_1022; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1024 = 4'hc == _T_88553 ? shiftedStoreDataKnownPReg_12 : _GEN_1023; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1025 = 4'hd == _T_88553 ? shiftedStoreDataKnownPReg_13 : _GEN_1024; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1026 = 4'he == _T_88553 ? shiftedStoreDataKnownPReg_14 : _GEN_1025; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1027 = 4'hf == _T_88553 ? shiftedStoreDataKnownPReg_15 : _GEN_1026; // @[LoadQueue.scala 194:31:@35349.6]
  assign _GEN_1029 = 4'h1 == _T_88553 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1030 = 4'h2 == _T_88553 ? shiftedStoreDataQPreg_2 : _GEN_1029; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1031 = 4'h3 == _T_88553 ? shiftedStoreDataQPreg_3 : _GEN_1030; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1032 = 4'h4 == _T_88553 ? shiftedStoreDataQPreg_4 : _GEN_1031; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1033 = 4'h5 == _T_88553 ? shiftedStoreDataQPreg_5 : _GEN_1032; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1034 = 4'h6 == _T_88553 ? shiftedStoreDataQPreg_6 : _GEN_1033; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1035 = 4'h7 == _T_88553 ? shiftedStoreDataQPreg_7 : _GEN_1034; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1036 = 4'h8 == _T_88553 ? shiftedStoreDataQPreg_8 : _GEN_1035; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1037 = 4'h9 == _T_88553 ? shiftedStoreDataQPreg_9 : _GEN_1036; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1038 = 4'ha == _T_88553 ? shiftedStoreDataQPreg_10 : _GEN_1037; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1039 = 4'hb == _T_88553 ? shiftedStoreDataQPreg_11 : _GEN_1038; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1040 = 4'hc == _T_88553 ? shiftedStoreDataQPreg_12 : _GEN_1039; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1041 = 4'hd == _T_88553 ? shiftedStoreDataQPreg_13 : _GEN_1040; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1042 = 4'he == _T_88553 ? shiftedStoreDataQPreg_14 : _GEN_1041; // @[LoadQueue.scala 195:31:@35350.6]
  assign _GEN_1043 = 4'hf == _T_88553 ? shiftedStoreDataQPreg_15 : _GEN_1042; // @[LoadQueue.scala 195:31:@35350.6]
  assign lastConflict_2_0 = _T_88570 ? _GEN_996 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_1 = _T_88570 ? _GEN_997 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_2 = _T_88570 ? _GEN_998 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_3 = _T_88570 ? _GEN_999 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_4 = _T_88570 ? _GEN_1000 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_5 = _T_88570 ? _GEN_1001 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_6 = _T_88570 ? _GEN_1002 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_7 = _T_88570 ? _GEN_1003 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_8 = _T_88570 ? _GEN_1004 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_9 = _T_88570 ? _GEN_1005 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_10 = _T_88570 ? _GEN_1006 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_11 = _T_88570 ? _GEN_1007 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_12 = _T_88570 ? _GEN_1008 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_13 = _T_88570 ? _GEN_1009 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_14 = _T_88570 ? _GEN_1010 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign lastConflict_2_15 = _T_88570 ? _GEN_1011 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign canBypass_2 = _T_88570 ? _GEN_1027 : 1'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign bypassVal_2 = _T_88570 ? _GEN_1043 : 32'h0; // @[LoadQueue.scala 192:53:@35347.4]
  assign _T_88676 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[LoadQueue.scala 191:60:@35404.4]
  assign _T_88677 = conflictPReg_3_3 ? 2'h3 : _T_88676; // @[LoadQueue.scala 191:60:@35405.4]
  assign _T_88678 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_88677}; // @[LoadQueue.scala 191:60:@35406.4]
  assign _T_88679 = conflictPReg_3_5 ? 3'h5 : _T_88678; // @[LoadQueue.scala 191:60:@35407.4]
  assign _T_88680 = conflictPReg_3_6 ? 3'h6 : _T_88679; // @[LoadQueue.scala 191:60:@35408.4]
  assign _T_88681 = conflictPReg_3_7 ? 3'h7 : _T_88680; // @[LoadQueue.scala 191:60:@35409.4]
  assign _T_88682 = conflictPReg_3_8 ? 4'h8 : {{1'd0}, _T_88681}; // @[LoadQueue.scala 191:60:@35410.4]
  assign _T_88683 = conflictPReg_3_9 ? 4'h9 : _T_88682; // @[LoadQueue.scala 191:60:@35411.4]
  assign _T_88684 = conflictPReg_3_10 ? 4'ha : _T_88683; // @[LoadQueue.scala 191:60:@35412.4]
  assign _T_88685 = conflictPReg_3_11 ? 4'hb : _T_88684; // @[LoadQueue.scala 191:60:@35413.4]
  assign _T_88686 = conflictPReg_3_12 ? 4'hc : _T_88685; // @[LoadQueue.scala 191:60:@35414.4]
  assign _T_88687 = conflictPReg_3_13 ? 4'hd : _T_88686; // @[LoadQueue.scala 191:60:@35415.4]
  assign _T_88688 = conflictPReg_3_14 ? 4'he : _T_88687; // @[LoadQueue.scala 191:60:@35416.4]
  assign _T_88689 = conflictPReg_3_15 ? 4'hf : _T_88688; // @[LoadQueue.scala 191:60:@35417.4]
  assign _T_88692 = conflictPReg_3_0 | conflictPReg_3_1; // @[LoadQueue.scala 192:43:@35419.4]
  assign _T_88693 = _T_88692 | conflictPReg_3_2; // @[LoadQueue.scala 192:43:@35420.4]
  assign _T_88694 = _T_88693 | conflictPReg_3_3; // @[LoadQueue.scala 192:43:@35421.4]
  assign _T_88695 = _T_88694 | conflictPReg_3_4; // @[LoadQueue.scala 192:43:@35422.4]
  assign _T_88696 = _T_88695 | conflictPReg_3_5; // @[LoadQueue.scala 192:43:@35423.4]
  assign _T_88697 = _T_88696 | conflictPReg_3_6; // @[LoadQueue.scala 192:43:@35424.4]
  assign _T_88698 = _T_88697 | conflictPReg_3_7; // @[LoadQueue.scala 192:43:@35425.4]
  assign _T_88699 = _T_88698 | conflictPReg_3_8; // @[LoadQueue.scala 192:43:@35426.4]
  assign _T_88700 = _T_88699 | conflictPReg_3_9; // @[LoadQueue.scala 192:43:@35427.4]
  assign _T_88701 = _T_88700 | conflictPReg_3_10; // @[LoadQueue.scala 192:43:@35428.4]
  assign _T_88702 = _T_88701 | conflictPReg_3_11; // @[LoadQueue.scala 192:43:@35429.4]
  assign _T_88703 = _T_88702 | conflictPReg_3_12; // @[LoadQueue.scala 192:43:@35430.4]
  assign _T_88704 = _T_88703 | conflictPReg_3_13; // @[LoadQueue.scala 192:43:@35431.4]
  assign _T_88705 = _T_88704 | conflictPReg_3_14; // @[LoadQueue.scala 192:43:@35432.4]
  assign _T_88706 = _T_88705 | conflictPReg_3_15; // @[LoadQueue.scala 192:43:@35433.4]
  assign _GEN_1062 = 4'h0 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1063 = 4'h1 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1064 = 4'h2 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1065 = 4'h3 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1066 = 4'h4 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1067 = 4'h5 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1068 = 4'h6 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1069 = 4'h7 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1070 = 4'h8 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1071 = 4'h9 == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1072 = 4'ha == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1073 = 4'hb == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1074 = 4'hc == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1075 = 4'hd == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1076 = 4'he == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1077 = 4'hf == _T_88689; // @[LoadQueue.scala 193:43:@35435.6]
  assign _GEN_1079 = 4'h1 == _T_88689 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1080 = 4'h2 == _T_88689 ? shiftedStoreDataKnownPReg_2 : _GEN_1079; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1081 = 4'h3 == _T_88689 ? shiftedStoreDataKnownPReg_3 : _GEN_1080; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1082 = 4'h4 == _T_88689 ? shiftedStoreDataKnownPReg_4 : _GEN_1081; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1083 = 4'h5 == _T_88689 ? shiftedStoreDataKnownPReg_5 : _GEN_1082; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1084 = 4'h6 == _T_88689 ? shiftedStoreDataKnownPReg_6 : _GEN_1083; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1085 = 4'h7 == _T_88689 ? shiftedStoreDataKnownPReg_7 : _GEN_1084; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1086 = 4'h8 == _T_88689 ? shiftedStoreDataKnownPReg_8 : _GEN_1085; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1087 = 4'h9 == _T_88689 ? shiftedStoreDataKnownPReg_9 : _GEN_1086; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1088 = 4'ha == _T_88689 ? shiftedStoreDataKnownPReg_10 : _GEN_1087; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1089 = 4'hb == _T_88689 ? shiftedStoreDataKnownPReg_11 : _GEN_1088; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1090 = 4'hc == _T_88689 ? shiftedStoreDataKnownPReg_12 : _GEN_1089; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1091 = 4'hd == _T_88689 ? shiftedStoreDataKnownPReg_13 : _GEN_1090; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1092 = 4'he == _T_88689 ? shiftedStoreDataKnownPReg_14 : _GEN_1091; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1093 = 4'hf == _T_88689 ? shiftedStoreDataKnownPReg_15 : _GEN_1092; // @[LoadQueue.scala 194:31:@35436.6]
  assign _GEN_1095 = 4'h1 == _T_88689 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1096 = 4'h2 == _T_88689 ? shiftedStoreDataQPreg_2 : _GEN_1095; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1097 = 4'h3 == _T_88689 ? shiftedStoreDataQPreg_3 : _GEN_1096; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1098 = 4'h4 == _T_88689 ? shiftedStoreDataQPreg_4 : _GEN_1097; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1099 = 4'h5 == _T_88689 ? shiftedStoreDataQPreg_5 : _GEN_1098; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1100 = 4'h6 == _T_88689 ? shiftedStoreDataQPreg_6 : _GEN_1099; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1101 = 4'h7 == _T_88689 ? shiftedStoreDataQPreg_7 : _GEN_1100; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1102 = 4'h8 == _T_88689 ? shiftedStoreDataQPreg_8 : _GEN_1101; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1103 = 4'h9 == _T_88689 ? shiftedStoreDataQPreg_9 : _GEN_1102; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1104 = 4'ha == _T_88689 ? shiftedStoreDataQPreg_10 : _GEN_1103; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1105 = 4'hb == _T_88689 ? shiftedStoreDataQPreg_11 : _GEN_1104; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1106 = 4'hc == _T_88689 ? shiftedStoreDataQPreg_12 : _GEN_1105; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1107 = 4'hd == _T_88689 ? shiftedStoreDataQPreg_13 : _GEN_1106; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1108 = 4'he == _T_88689 ? shiftedStoreDataQPreg_14 : _GEN_1107; // @[LoadQueue.scala 195:31:@35437.6]
  assign _GEN_1109 = 4'hf == _T_88689 ? shiftedStoreDataQPreg_15 : _GEN_1108; // @[LoadQueue.scala 195:31:@35437.6]
  assign lastConflict_3_0 = _T_88706 ? _GEN_1062 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_1 = _T_88706 ? _GEN_1063 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_2 = _T_88706 ? _GEN_1064 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_3 = _T_88706 ? _GEN_1065 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_4 = _T_88706 ? _GEN_1066 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_5 = _T_88706 ? _GEN_1067 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_6 = _T_88706 ? _GEN_1068 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_7 = _T_88706 ? _GEN_1069 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_8 = _T_88706 ? _GEN_1070 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_9 = _T_88706 ? _GEN_1071 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_10 = _T_88706 ? _GEN_1072 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_11 = _T_88706 ? _GEN_1073 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_12 = _T_88706 ? _GEN_1074 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_13 = _T_88706 ? _GEN_1075 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_14 = _T_88706 ? _GEN_1076 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign lastConflict_3_15 = _T_88706 ? _GEN_1077 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign canBypass_3 = _T_88706 ? _GEN_1093 : 1'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign bypassVal_3 = _T_88706 ? _GEN_1109 : 32'h0; // @[LoadQueue.scala 192:53:@35434.4]
  assign _T_88812 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[LoadQueue.scala 191:60:@35491.4]
  assign _T_88813 = conflictPReg_4_3 ? 2'h3 : _T_88812; // @[LoadQueue.scala 191:60:@35492.4]
  assign _T_88814 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_88813}; // @[LoadQueue.scala 191:60:@35493.4]
  assign _T_88815 = conflictPReg_4_5 ? 3'h5 : _T_88814; // @[LoadQueue.scala 191:60:@35494.4]
  assign _T_88816 = conflictPReg_4_6 ? 3'h6 : _T_88815; // @[LoadQueue.scala 191:60:@35495.4]
  assign _T_88817 = conflictPReg_4_7 ? 3'h7 : _T_88816; // @[LoadQueue.scala 191:60:@35496.4]
  assign _T_88818 = conflictPReg_4_8 ? 4'h8 : {{1'd0}, _T_88817}; // @[LoadQueue.scala 191:60:@35497.4]
  assign _T_88819 = conflictPReg_4_9 ? 4'h9 : _T_88818; // @[LoadQueue.scala 191:60:@35498.4]
  assign _T_88820 = conflictPReg_4_10 ? 4'ha : _T_88819; // @[LoadQueue.scala 191:60:@35499.4]
  assign _T_88821 = conflictPReg_4_11 ? 4'hb : _T_88820; // @[LoadQueue.scala 191:60:@35500.4]
  assign _T_88822 = conflictPReg_4_12 ? 4'hc : _T_88821; // @[LoadQueue.scala 191:60:@35501.4]
  assign _T_88823 = conflictPReg_4_13 ? 4'hd : _T_88822; // @[LoadQueue.scala 191:60:@35502.4]
  assign _T_88824 = conflictPReg_4_14 ? 4'he : _T_88823; // @[LoadQueue.scala 191:60:@35503.4]
  assign _T_88825 = conflictPReg_4_15 ? 4'hf : _T_88824; // @[LoadQueue.scala 191:60:@35504.4]
  assign _T_88828 = conflictPReg_4_0 | conflictPReg_4_1; // @[LoadQueue.scala 192:43:@35506.4]
  assign _T_88829 = _T_88828 | conflictPReg_4_2; // @[LoadQueue.scala 192:43:@35507.4]
  assign _T_88830 = _T_88829 | conflictPReg_4_3; // @[LoadQueue.scala 192:43:@35508.4]
  assign _T_88831 = _T_88830 | conflictPReg_4_4; // @[LoadQueue.scala 192:43:@35509.4]
  assign _T_88832 = _T_88831 | conflictPReg_4_5; // @[LoadQueue.scala 192:43:@35510.4]
  assign _T_88833 = _T_88832 | conflictPReg_4_6; // @[LoadQueue.scala 192:43:@35511.4]
  assign _T_88834 = _T_88833 | conflictPReg_4_7; // @[LoadQueue.scala 192:43:@35512.4]
  assign _T_88835 = _T_88834 | conflictPReg_4_8; // @[LoadQueue.scala 192:43:@35513.4]
  assign _T_88836 = _T_88835 | conflictPReg_4_9; // @[LoadQueue.scala 192:43:@35514.4]
  assign _T_88837 = _T_88836 | conflictPReg_4_10; // @[LoadQueue.scala 192:43:@35515.4]
  assign _T_88838 = _T_88837 | conflictPReg_4_11; // @[LoadQueue.scala 192:43:@35516.4]
  assign _T_88839 = _T_88838 | conflictPReg_4_12; // @[LoadQueue.scala 192:43:@35517.4]
  assign _T_88840 = _T_88839 | conflictPReg_4_13; // @[LoadQueue.scala 192:43:@35518.4]
  assign _T_88841 = _T_88840 | conflictPReg_4_14; // @[LoadQueue.scala 192:43:@35519.4]
  assign _T_88842 = _T_88841 | conflictPReg_4_15; // @[LoadQueue.scala 192:43:@35520.4]
  assign _GEN_1128 = 4'h0 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1129 = 4'h1 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1130 = 4'h2 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1131 = 4'h3 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1132 = 4'h4 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1133 = 4'h5 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1134 = 4'h6 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1135 = 4'h7 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1136 = 4'h8 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1137 = 4'h9 == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1138 = 4'ha == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1139 = 4'hb == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1140 = 4'hc == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1141 = 4'hd == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1142 = 4'he == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1143 = 4'hf == _T_88825; // @[LoadQueue.scala 193:43:@35522.6]
  assign _GEN_1145 = 4'h1 == _T_88825 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1146 = 4'h2 == _T_88825 ? shiftedStoreDataKnownPReg_2 : _GEN_1145; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1147 = 4'h3 == _T_88825 ? shiftedStoreDataKnownPReg_3 : _GEN_1146; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1148 = 4'h4 == _T_88825 ? shiftedStoreDataKnownPReg_4 : _GEN_1147; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1149 = 4'h5 == _T_88825 ? shiftedStoreDataKnownPReg_5 : _GEN_1148; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1150 = 4'h6 == _T_88825 ? shiftedStoreDataKnownPReg_6 : _GEN_1149; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1151 = 4'h7 == _T_88825 ? shiftedStoreDataKnownPReg_7 : _GEN_1150; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1152 = 4'h8 == _T_88825 ? shiftedStoreDataKnownPReg_8 : _GEN_1151; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1153 = 4'h9 == _T_88825 ? shiftedStoreDataKnownPReg_9 : _GEN_1152; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1154 = 4'ha == _T_88825 ? shiftedStoreDataKnownPReg_10 : _GEN_1153; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1155 = 4'hb == _T_88825 ? shiftedStoreDataKnownPReg_11 : _GEN_1154; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1156 = 4'hc == _T_88825 ? shiftedStoreDataKnownPReg_12 : _GEN_1155; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1157 = 4'hd == _T_88825 ? shiftedStoreDataKnownPReg_13 : _GEN_1156; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1158 = 4'he == _T_88825 ? shiftedStoreDataKnownPReg_14 : _GEN_1157; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1159 = 4'hf == _T_88825 ? shiftedStoreDataKnownPReg_15 : _GEN_1158; // @[LoadQueue.scala 194:31:@35523.6]
  assign _GEN_1161 = 4'h1 == _T_88825 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1162 = 4'h2 == _T_88825 ? shiftedStoreDataQPreg_2 : _GEN_1161; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1163 = 4'h3 == _T_88825 ? shiftedStoreDataQPreg_3 : _GEN_1162; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1164 = 4'h4 == _T_88825 ? shiftedStoreDataQPreg_4 : _GEN_1163; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1165 = 4'h5 == _T_88825 ? shiftedStoreDataQPreg_5 : _GEN_1164; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1166 = 4'h6 == _T_88825 ? shiftedStoreDataQPreg_6 : _GEN_1165; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1167 = 4'h7 == _T_88825 ? shiftedStoreDataQPreg_7 : _GEN_1166; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1168 = 4'h8 == _T_88825 ? shiftedStoreDataQPreg_8 : _GEN_1167; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1169 = 4'h9 == _T_88825 ? shiftedStoreDataQPreg_9 : _GEN_1168; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1170 = 4'ha == _T_88825 ? shiftedStoreDataQPreg_10 : _GEN_1169; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1171 = 4'hb == _T_88825 ? shiftedStoreDataQPreg_11 : _GEN_1170; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1172 = 4'hc == _T_88825 ? shiftedStoreDataQPreg_12 : _GEN_1171; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1173 = 4'hd == _T_88825 ? shiftedStoreDataQPreg_13 : _GEN_1172; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1174 = 4'he == _T_88825 ? shiftedStoreDataQPreg_14 : _GEN_1173; // @[LoadQueue.scala 195:31:@35524.6]
  assign _GEN_1175 = 4'hf == _T_88825 ? shiftedStoreDataQPreg_15 : _GEN_1174; // @[LoadQueue.scala 195:31:@35524.6]
  assign lastConflict_4_0 = _T_88842 ? _GEN_1128 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_1 = _T_88842 ? _GEN_1129 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_2 = _T_88842 ? _GEN_1130 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_3 = _T_88842 ? _GEN_1131 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_4 = _T_88842 ? _GEN_1132 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_5 = _T_88842 ? _GEN_1133 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_6 = _T_88842 ? _GEN_1134 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_7 = _T_88842 ? _GEN_1135 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_8 = _T_88842 ? _GEN_1136 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_9 = _T_88842 ? _GEN_1137 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_10 = _T_88842 ? _GEN_1138 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_11 = _T_88842 ? _GEN_1139 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_12 = _T_88842 ? _GEN_1140 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_13 = _T_88842 ? _GEN_1141 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_14 = _T_88842 ? _GEN_1142 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign lastConflict_4_15 = _T_88842 ? _GEN_1143 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign canBypass_4 = _T_88842 ? _GEN_1159 : 1'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign bypassVal_4 = _T_88842 ? _GEN_1175 : 32'h0; // @[LoadQueue.scala 192:53:@35521.4]
  assign _T_88948 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[LoadQueue.scala 191:60:@35578.4]
  assign _T_88949 = conflictPReg_5_3 ? 2'h3 : _T_88948; // @[LoadQueue.scala 191:60:@35579.4]
  assign _T_88950 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_88949}; // @[LoadQueue.scala 191:60:@35580.4]
  assign _T_88951 = conflictPReg_5_5 ? 3'h5 : _T_88950; // @[LoadQueue.scala 191:60:@35581.4]
  assign _T_88952 = conflictPReg_5_6 ? 3'h6 : _T_88951; // @[LoadQueue.scala 191:60:@35582.4]
  assign _T_88953 = conflictPReg_5_7 ? 3'h7 : _T_88952; // @[LoadQueue.scala 191:60:@35583.4]
  assign _T_88954 = conflictPReg_5_8 ? 4'h8 : {{1'd0}, _T_88953}; // @[LoadQueue.scala 191:60:@35584.4]
  assign _T_88955 = conflictPReg_5_9 ? 4'h9 : _T_88954; // @[LoadQueue.scala 191:60:@35585.4]
  assign _T_88956 = conflictPReg_5_10 ? 4'ha : _T_88955; // @[LoadQueue.scala 191:60:@35586.4]
  assign _T_88957 = conflictPReg_5_11 ? 4'hb : _T_88956; // @[LoadQueue.scala 191:60:@35587.4]
  assign _T_88958 = conflictPReg_5_12 ? 4'hc : _T_88957; // @[LoadQueue.scala 191:60:@35588.4]
  assign _T_88959 = conflictPReg_5_13 ? 4'hd : _T_88958; // @[LoadQueue.scala 191:60:@35589.4]
  assign _T_88960 = conflictPReg_5_14 ? 4'he : _T_88959; // @[LoadQueue.scala 191:60:@35590.4]
  assign _T_88961 = conflictPReg_5_15 ? 4'hf : _T_88960; // @[LoadQueue.scala 191:60:@35591.4]
  assign _T_88964 = conflictPReg_5_0 | conflictPReg_5_1; // @[LoadQueue.scala 192:43:@35593.4]
  assign _T_88965 = _T_88964 | conflictPReg_5_2; // @[LoadQueue.scala 192:43:@35594.4]
  assign _T_88966 = _T_88965 | conflictPReg_5_3; // @[LoadQueue.scala 192:43:@35595.4]
  assign _T_88967 = _T_88966 | conflictPReg_5_4; // @[LoadQueue.scala 192:43:@35596.4]
  assign _T_88968 = _T_88967 | conflictPReg_5_5; // @[LoadQueue.scala 192:43:@35597.4]
  assign _T_88969 = _T_88968 | conflictPReg_5_6; // @[LoadQueue.scala 192:43:@35598.4]
  assign _T_88970 = _T_88969 | conflictPReg_5_7; // @[LoadQueue.scala 192:43:@35599.4]
  assign _T_88971 = _T_88970 | conflictPReg_5_8; // @[LoadQueue.scala 192:43:@35600.4]
  assign _T_88972 = _T_88971 | conflictPReg_5_9; // @[LoadQueue.scala 192:43:@35601.4]
  assign _T_88973 = _T_88972 | conflictPReg_5_10; // @[LoadQueue.scala 192:43:@35602.4]
  assign _T_88974 = _T_88973 | conflictPReg_5_11; // @[LoadQueue.scala 192:43:@35603.4]
  assign _T_88975 = _T_88974 | conflictPReg_5_12; // @[LoadQueue.scala 192:43:@35604.4]
  assign _T_88976 = _T_88975 | conflictPReg_5_13; // @[LoadQueue.scala 192:43:@35605.4]
  assign _T_88977 = _T_88976 | conflictPReg_5_14; // @[LoadQueue.scala 192:43:@35606.4]
  assign _T_88978 = _T_88977 | conflictPReg_5_15; // @[LoadQueue.scala 192:43:@35607.4]
  assign _GEN_1194 = 4'h0 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1195 = 4'h1 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1196 = 4'h2 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1197 = 4'h3 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1198 = 4'h4 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1199 = 4'h5 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1200 = 4'h6 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1201 = 4'h7 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1202 = 4'h8 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1203 = 4'h9 == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1204 = 4'ha == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1205 = 4'hb == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1206 = 4'hc == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1207 = 4'hd == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1208 = 4'he == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1209 = 4'hf == _T_88961; // @[LoadQueue.scala 193:43:@35609.6]
  assign _GEN_1211 = 4'h1 == _T_88961 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1212 = 4'h2 == _T_88961 ? shiftedStoreDataKnownPReg_2 : _GEN_1211; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1213 = 4'h3 == _T_88961 ? shiftedStoreDataKnownPReg_3 : _GEN_1212; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1214 = 4'h4 == _T_88961 ? shiftedStoreDataKnownPReg_4 : _GEN_1213; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1215 = 4'h5 == _T_88961 ? shiftedStoreDataKnownPReg_5 : _GEN_1214; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1216 = 4'h6 == _T_88961 ? shiftedStoreDataKnownPReg_6 : _GEN_1215; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1217 = 4'h7 == _T_88961 ? shiftedStoreDataKnownPReg_7 : _GEN_1216; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1218 = 4'h8 == _T_88961 ? shiftedStoreDataKnownPReg_8 : _GEN_1217; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1219 = 4'h9 == _T_88961 ? shiftedStoreDataKnownPReg_9 : _GEN_1218; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1220 = 4'ha == _T_88961 ? shiftedStoreDataKnownPReg_10 : _GEN_1219; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1221 = 4'hb == _T_88961 ? shiftedStoreDataKnownPReg_11 : _GEN_1220; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1222 = 4'hc == _T_88961 ? shiftedStoreDataKnownPReg_12 : _GEN_1221; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1223 = 4'hd == _T_88961 ? shiftedStoreDataKnownPReg_13 : _GEN_1222; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1224 = 4'he == _T_88961 ? shiftedStoreDataKnownPReg_14 : _GEN_1223; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1225 = 4'hf == _T_88961 ? shiftedStoreDataKnownPReg_15 : _GEN_1224; // @[LoadQueue.scala 194:31:@35610.6]
  assign _GEN_1227 = 4'h1 == _T_88961 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1228 = 4'h2 == _T_88961 ? shiftedStoreDataQPreg_2 : _GEN_1227; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1229 = 4'h3 == _T_88961 ? shiftedStoreDataQPreg_3 : _GEN_1228; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1230 = 4'h4 == _T_88961 ? shiftedStoreDataQPreg_4 : _GEN_1229; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1231 = 4'h5 == _T_88961 ? shiftedStoreDataQPreg_5 : _GEN_1230; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1232 = 4'h6 == _T_88961 ? shiftedStoreDataQPreg_6 : _GEN_1231; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1233 = 4'h7 == _T_88961 ? shiftedStoreDataQPreg_7 : _GEN_1232; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1234 = 4'h8 == _T_88961 ? shiftedStoreDataQPreg_8 : _GEN_1233; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1235 = 4'h9 == _T_88961 ? shiftedStoreDataQPreg_9 : _GEN_1234; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1236 = 4'ha == _T_88961 ? shiftedStoreDataQPreg_10 : _GEN_1235; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1237 = 4'hb == _T_88961 ? shiftedStoreDataQPreg_11 : _GEN_1236; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1238 = 4'hc == _T_88961 ? shiftedStoreDataQPreg_12 : _GEN_1237; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1239 = 4'hd == _T_88961 ? shiftedStoreDataQPreg_13 : _GEN_1238; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1240 = 4'he == _T_88961 ? shiftedStoreDataQPreg_14 : _GEN_1239; // @[LoadQueue.scala 195:31:@35611.6]
  assign _GEN_1241 = 4'hf == _T_88961 ? shiftedStoreDataQPreg_15 : _GEN_1240; // @[LoadQueue.scala 195:31:@35611.6]
  assign lastConflict_5_0 = _T_88978 ? _GEN_1194 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_1 = _T_88978 ? _GEN_1195 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_2 = _T_88978 ? _GEN_1196 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_3 = _T_88978 ? _GEN_1197 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_4 = _T_88978 ? _GEN_1198 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_5 = _T_88978 ? _GEN_1199 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_6 = _T_88978 ? _GEN_1200 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_7 = _T_88978 ? _GEN_1201 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_8 = _T_88978 ? _GEN_1202 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_9 = _T_88978 ? _GEN_1203 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_10 = _T_88978 ? _GEN_1204 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_11 = _T_88978 ? _GEN_1205 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_12 = _T_88978 ? _GEN_1206 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_13 = _T_88978 ? _GEN_1207 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_14 = _T_88978 ? _GEN_1208 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign lastConflict_5_15 = _T_88978 ? _GEN_1209 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign canBypass_5 = _T_88978 ? _GEN_1225 : 1'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign bypassVal_5 = _T_88978 ? _GEN_1241 : 32'h0; // @[LoadQueue.scala 192:53:@35608.4]
  assign _T_89084 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[LoadQueue.scala 191:60:@35665.4]
  assign _T_89085 = conflictPReg_6_3 ? 2'h3 : _T_89084; // @[LoadQueue.scala 191:60:@35666.4]
  assign _T_89086 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_89085}; // @[LoadQueue.scala 191:60:@35667.4]
  assign _T_89087 = conflictPReg_6_5 ? 3'h5 : _T_89086; // @[LoadQueue.scala 191:60:@35668.4]
  assign _T_89088 = conflictPReg_6_6 ? 3'h6 : _T_89087; // @[LoadQueue.scala 191:60:@35669.4]
  assign _T_89089 = conflictPReg_6_7 ? 3'h7 : _T_89088; // @[LoadQueue.scala 191:60:@35670.4]
  assign _T_89090 = conflictPReg_6_8 ? 4'h8 : {{1'd0}, _T_89089}; // @[LoadQueue.scala 191:60:@35671.4]
  assign _T_89091 = conflictPReg_6_9 ? 4'h9 : _T_89090; // @[LoadQueue.scala 191:60:@35672.4]
  assign _T_89092 = conflictPReg_6_10 ? 4'ha : _T_89091; // @[LoadQueue.scala 191:60:@35673.4]
  assign _T_89093 = conflictPReg_6_11 ? 4'hb : _T_89092; // @[LoadQueue.scala 191:60:@35674.4]
  assign _T_89094 = conflictPReg_6_12 ? 4'hc : _T_89093; // @[LoadQueue.scala 191:60:@35675.4]
  assign _T_89095 = conflictPReg_6_13 ? 4'hd : _T_89094; // @[LoadQueue.scala 191:60:@35676.4]
  assign _T_89096 = conflictPReg_6_14 ? 4'he : _T_89095; // @[LoadQueue.scala 191:60:@35677.4]
  assign _T_89097 = conflictPReg_6_15 ? 4'hf : _T_89096; // @[LoadQueue.scala 191:60:@35678.4]
  assign _T_89100 = conflictPReg_6_0 | conflictPReg_6_1; // @[LoadQueue.scala 192:43:@35680.4]
  assign _T_89101 = _T_89100 | conflictPReg_6_2; // @[LoadQueue.scala 192:43:@35681.4]
  assign _T_89102 = _T_89101 | conflictPReg_6_3; // @[LoadQueue.scala 192:43:@35682.4]
  assign _T_89103 = _T_89102 | conflictPReg_6_4; // @[LoadQueue.scala 192:43:@35683.4]
  assign _T_89104 = _T_89103 | conflictPReg_6_5; // @[LoadQueue.scala 192:43:@35684.4]
  assign _T_89105 = _T_89104 | conflictPReg_6_6; // @[LoadQueue.scala 192:43:@35685.4]
  assign _T_89106 = _T_89105 | conflictPReg_6_7; // @[LoadQueue.scala 192:43:@35686.4]
  assign _T_89107 = _T_89106 | conflictPReg_6_8; // @[LoadQueue.scala 192:43:@35687.4]
  assign _T_89108 = _T_89107 | conflictPReg_6_9; // @[LoadQueue.scala 192:43:@35688.4]
  assign _T_89109 = _T_89108 | conflictPReg_6_10; // @[LoadQueue.scala 192:43:@35689.4]
  assign _T_89110 = _T_89109 | conflictPReg_6_11; // @[LoadQueue.scala 192:43:@35690.4]
  assign _T_89111 = _T_89110 | conflictPReg_6_12; // @[LoadQueue.scala 192:43:@35691.4]
  assign _T_89112 = _T_89111 | conflictPReg_6_13; // @[LoadQueue.scala 192:43:@35692.4]
  assign _T_89113 = _T_89112 | conflictPReg_6_14; // @[LoadQueue.scala 192:43:@35693.4]
  assign _T_89114 = _T_89113 | conflictPReg_6_15; // @[LoadQueue.scala 192:43:@35694.4]
  assign _GEN_1260 = 4'h0 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1261 = 4'h1 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1262 = 4'h2 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1263 = 4'h3 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1264 = 4'h4 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1265 = 4'h5 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1266 = 4'h6 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1267 = 4'h7 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1268 = 4'h8 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1269 = 4'h9 == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1270 = 4'ha == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1271 = 4'hb == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1272 = 4'hc == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1273 = 4'hd == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1274 = 4'he == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1275 = 4'hf == _T_89097; // @[LoadQueue.scala 193:43:@35696.6]
  assign _GEN_1277 = 4'h1 == _T_89097 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1278 = 4'h2 == _T_89097 ? shiftedStoreDataKnownPReg_2 : _GEN_1277; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1279 = 4'h3 == _T_89097 ? shiftedStoreDataKnownPReg_3 : _GEN_1278; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1280 = 4'h4 == _T_89097 ? shiftedStoreDataKnownPReg_4 : _GEN_1279; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1281 = 4'h5 == _T_89097 ? shiftedStoreDataKnownPReg_5 : _GEN_1280; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1282 = 4'h6 == _T_89097 ? shiftedStoreDataKnownPReg_6 : _GEN_1281; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1283 = 4'h7 == _T_89097 ? shiftedStoreDataKnownPReg_7 : _GEN_1282; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1284 = 4'h8 == _T_89097 ? shiftedStoreDataKnownPReg_8 : _GEN_1283; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1285 = 4'h9 == _T_89097 ? shiftedStoreDataKnownPReg_9 : _GEN_1284; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1286 = 4'ha == _T_89097 ? shiftedStoreDataKnownPReg_10 : _GEN_1285; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1287 = 4'hb == _T_89097 ? shiftedStoreDataKnownPReg_11 : _GEN_1286; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1288 = 4'hc == _T_89097 ? shiftedStoreDataKnownPReg_12 : _GEN_1287; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1289 = 4'hd == _T_89097 ? shiftedStoreDataKnownPReg_13 : _GEN_1288; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1290 = 4'he == _T_89097 ? shiftedStoreDataKnownPReg_14 : _GEN_1289; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1291 = 4'hf == _T_89097 ? shiftedStoreDataKnownPReg_15 : _GEN_1290; // @[LoadQueue.scala 194:31:@35697.6]
  assign _GEN_1293 = 4'h1 == _T_89097 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1294 = 4'h2 == _T_89097 ? shiftedStoreDataQPreg_2 : _GEN_1293; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1295 = 4'h3 == _T_89097 ? shiftedStoreDataQPreg_3 : _GEN_1294; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1296 = 4'h4 == _T_89097 ? shiftedStoreDataQPreg_4 : _GEN_1295; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1297 = 4'h5 == _T_89097 ? shiftedStoreDataQPreg_5 : _GEN_1296; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1298 = 4'h6 == _T_89097 ? shiftedStoreDataQPreg_6 : _GEN_1297; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1299 = 4'h7 == _T_89097 ? shiftedStoreDataQPreg_7 : _GEN_1298; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1300 = 4'h8 == _T_89097 ? shiftedStoreDataQPreg_8 : _GEN_1299; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1301 = 4'h9 == _T_89097 ? shiftedStoreDataQPreg_9 : _GEN_1300; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1302 = 4'ha == _T_89097 ? shiftedStoreDataQPreg_10 : _GEN_1301; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1303 = 4'hb == _T_89097 ? shiftedStoreDataQPreg_11 : _GEN_1302; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1304 = 4'hc == _T_89097 ? shiftedStoreDataQPreg_12 : _GEN_1303; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1305 = 4'hd == _T_89097 ? shiftedStoreDataQPreg_13 : _GEN_1304; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1306 = 4'he == _T_89097 ? shiftedStoreDataQPreg_14 : _GEN_1305; // @[LoadQueue.scala 195:31:@35698.6]
  assign _GEN_1307 = 4'hf == _T_89097 ? shiftedStoreDataQPreg_15 : _GEN_1306; // @[LoadQueue.scala 195:31:@35698.6]
  assign lastConflict_6_0 = _T_89114 ? _GEN_1260 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_1 = _T_89114 ? _GEN_1261 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_2 = _T_89114 ? _GEN_1262 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_3 = _T_89114 ? _GEN_1263 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_4 = _T_89114 ? _GEN_1264 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_5 = _T_89114 ? _GEN_1265 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_6 = _T_89114 ? _GEN_1266 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_7 = _T_89114 ? _GEN_1267 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_8 = _T_89114 ? _GEN_1268 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_9 = _T_89114 ? _GEN_1269 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_10 = _T_89114 ? _GEN_1270 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_11 = _T_89114 ? _GEN_1271 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_12 = _T_89114 ? _GEN_1272 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_13 = _T_89114 ? _GEN_1273 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_14 = _T_89114 ? _GEN_1274 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign lastConflict_6_15 = _T_89114 ? _GEN_1275 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign canBypass_6 = _T_89114 ? _GEN_1291 : 1'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign bypassVal_6 = _T_89114 ? _GEN_1307 : 32'h0; // @[LoadQueue.scala 192:53:@35695.4]
  assign _T_89220 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[LoadQueue.scala 191:60:@35752.4]
  assign _T_89221 = conflictPReg_7_3 ? 2'h3 : _T_89220; // @[LoadQueue.scala 191:60:@35753.4]
  assign _T_89222 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_89221}; // @[LoadQueue.scala 191:60:@35754.4]
  assign _T_89223 = conflictPReg_7_5 ? 3'h5 : _T_89222; // @[LoadQueue.scala 191:60:@35755.4]
  assign _T_89224 = conflictPReg_7_6 ? 3'h6 : _T_89223; // @[LoadQueue.scala 191:60:@35756.4]
  assign _T_89225 = conflictPReg_7_7 ? 3'h7 : _T_89224; // @[LoadQueue.scala 191:60:@35757.4]
  assign _T_89226 = conflictPReg_7_8 ? 4'h8 : {{1'd0}, _T_89225}; // @[LoadQueue.scala 191:60:@35758.4]
  assign _T_89227 = conflictPReg_7_9 ? 4'h9 : _T_89226; // @[LoadQueue.scala 191:60:@35759.4]
  assign _T_89228 = conflictPReg_7_10 ? 4'ha : _T_89227; // @[LoadQueue.scala 191:60:@35760.4]
  assign _T_89229 = conflictPReg_7_11 ? 4'hb : _T_89228; // @[LoadQueue.scala 191:60:@35761.4]
  assign _T_89230 = conflictPReg_7_12 ? 4'hc : _T_89229; // @[LoadQueue.scala 191:60:@35762.4]
  assign _T_89231 = conflictPReg_7_13 ? 4'hd : _T_89230; // @[LoadQueue.scala 191:60:@35763.4]
  assign _T_89232 = conflictPReg_7_14 ? 4'he : _T_89231; // @[LoadQueue.scala 191:60:@35764.4]
  assign _T_89233 = conflictPReg_7_15 ? 4'hf : _T_89232; // @[LoadQueue.scala 191:60:@35765.4]
  assign _T_89236 = conflictPReg_7_0 | conflictPReg_7_1; // @[LoadQueue.scala 192:43:@35767.4]
  assign _T_89237 = _T_89236 | conflictPReg_7_2; // @[LoadQueue.scala 192:43:@35768.4]
  assign _T_89238 = _T_89237 | conflictPReg_7_3; // @[LoadQueue.scala 192:43:@35769.4]
  assign _T_89239 = _T_89238 | conflictPReg_7_4; // @[LoadQueue.scala 192:43:@35770.4]
  assign _T_89240 = _T_89239 | conflictPReg_7_5; // @[LoadQueue.scala 192:43:@35771.4]
  assign _T_89241 = _T_89240 | conflictPReg_7_6; // @[LoadQueue.scala 192:43:@35772.4]
  assign _T_89242 = _T_89241 | conflictPReg_7_7; // @[LoadQueue.scala 192:43:@35773.4]
  assign _T_89243 = _T_89242 | conflictPReg_7_8; // @[LoadQueue.scala 192:43:@35774.4]
  assign _T_89244 = _T_89243 | conflictPReg_7_9; // @[LoadQueue.scala 192:43:@35775.4]
  assign _T_89245 = _T_89244 | conflictPReg_7_10; // @[LoadQueue.scala 192:43:@35776.4]
  assign _T_89246 = _T_89245 | conflictPReg_7_11; // @[LoadQueue.scala 192:43:@35777.4]
  assign _T_89247 = _T_89246 | conflictPReg_7_12; // @[LoadQueue.scala 192:43:@35778.4]
  assign _T_89248 = _T_89247 | conflictPReg_7_13; // @[LoadQueue.scala 192:43:@35779.4]
  assign _T_89249 = _T_89248 | conflictPReg_7_14; // @[LoadQueue.scala 192:43:@35780.4]
  assign _T_89250 = _T_89249 | conflictPReg_7_15; // @[LoadQueue.scala 192:43:@35781.4]
  assign _GEN_1326 = 4'h0 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1327 = 4'h1 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1328 = 4'h2 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1329 = 4'h3 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1330 = 4'h4 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1331 = 4'h5 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1332 = 4'h6 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1333 = 4'h7 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1334 = 4'h8 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1335 = 4'h9 == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1336 = 4'ha == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1337 = 4'hb == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1338 = 4'hc == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1339 = 4'hd == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1340 = 4'he == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1341 = 4'hf == _T_89233; // @[LoadQueue.scala 193:43:@35783.6]
  assign _GEN_1343 = 4'h1 == _T_89233 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1344 = 4'h2 == _T_89233 ? shiftedStoreDataKnownPReg_2 : _GEN_1343; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1345 = 4'h3 == _T_89233 ? shiftedStoreDataKnownPReg_3 : _GEN_1344; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1346 = 4'h4 == _T_89233 ? shiftedStoreDataKnownPReg_4 : _GEN_1345; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1347 = 4'h5 == _T_89233 ? shiftedStoreDataKnownPReg_5 : _GEN_1346; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1348 = 4'h6 == _T_89233 ? shiftedStoreDataKnownPReg_6 : _GEN_1347; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1349 = 4'h7 == _T_89233 ? shiftedStoreDataKnownPReg_7 : _GEN_1348; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1350 = 4'h8 == _T_89233 ? shiftedStoreDataKnownPReg_8 : _GEN_1349; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1351 = 4'h9 == _T_89233 ? shiftedStoreDataKnownPReg_9 : _GEN_1350; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1352 = 4'ha == _T_89233 ? shiftedStoreDataKnownPReg_10 : _GEN_1351; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1353 = 4'hb == _T_89233 ? shiftedStoreDataKnownPReg_11 : _GEN_1352; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1354 = 4'hc == _T_89233 ? shiftedStoreDataKnownPReg_12 : _GEN_1353; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1355 = 4'hd == _T_89233 ? shiftedStoreDataKnownPReg_13 : _GEN_1354; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1356 = 4'he == _T_89233 ? shiftedStoreDataKnownPReg_14 : _GEN_1355; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1357 = 4'hf == _T_89233 ? shiftedStoreDataKnownPReg_15 : _GEN_1356; // @[LoadQueue.scala 194:31:@35784.6]
  assign _GEN_1359 = 4'h1 == _T_89233 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1360 = 4'h2 == _T_89233 ? shiftedStoreDataQPreg_2 : _GEN_1359; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1361 = 4'h3 == _T_89233 ? shiftedStoreDataQPreg_3 : _GEN_1360; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1362 = 4'h4 == _T_89233 ? shiftedStoreDataQPreg_4 : _GEN_1361; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1363 = 4'h5 == _T_89233 ? shiftedStoreDataQPreg_5 : _GEN_1362; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1364 = 4'h6 == _T_89233 ? shiftedStoreDataQPreg_6 : _GEN_1363; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1365 = 4'h7 == _T_89233 ? shiftedStoreDataQPreg_7 : _GEN_1364; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1366 = 4'h8 == _T_89233 ? shiftedStoreDataQPreg_8 : _GEN_1365; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1367 = 4'h9 == _T_89233 ? shiftedStoreDataQPreg_9 : _GEN_1366; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1368 = 4'ha == _T_89233 ? shiftedStoreDataQPreg_10 : _GEN_1367; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1369 = 4'hb == _T_89233 ? shiftedStoreDataQPreg_11 : _GEN_1368; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1370 = 4'hc == _T_89233 ? shiftedStoreDataQPreg_12 : _GEN_1369; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1371 = 4'hd == _T_89233 ? shiftedStoreDataQPreg_13 : _GEN_1370; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1372 = 4'he == _T_89233 ? shiftedStoreDataQPreg_14 : _GEN_1371; // @[LoadQueue.scala 195:31:@35785.6]
  assign _GEN_1373 = 4'hf == _T_89233 ? shiftedStoreDataQPreg_15 : _GEN_1372; // @[LoadQueue.scala 195:31:@35785.6]
  assign lastConflict_7_0 = _T_89250 ? _GEN_1326 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_1 = _T_89250 ? _GEN_1327 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_2 = _T_89250 ? _GEN_1328 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_3 = _T_89250 ? _GEN_1329 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_4 = _T_89250 ? _GEN_1330 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_5 = _T_89250 ? _GEN_1331 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_6 = _T_89250 ? _GEN_1332 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_7 = _T_89250 ? _GEN_1333 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_8 = _T_89250 ? _GEN_1334 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_9 = _T_89250 ? _GEN_1335 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_10 = _T_89250 ? _GEN_1336 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_11 = _T_89250 ? _GEN_1337 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_12 = _T_89250 ? _GEN_1338 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_13 = _T_89250 ? _GEN_1339 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_14 = _T_89250 ? _GEN_1340 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign lastConflict_7_15 = _T_89250 ? _GEN_1341 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign canBypass_7 = _T_89250 ? _GEN_1357 : 1'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign bypassVal_7 = _T_89250 ? _GEN_1373 : 32'h0; // @[LoadQueue.scala 192:53:@35782.4]
  assign _T_89356 = conflictPReg_8_2 ? 2'h2 : {{1'd0}, conflictPReg_8_1}; // @[LoadQueue.scala 191:60:@35839.4]
  assign _T_89357 = conflictPReg_8_3 ? 2'h3 : _T_89356; // @[LoadQueue.scala 191:60:@35840.4]
  assign _T_89358 = conflictPReg_8_4 ? 3'h4 : {{1'd0}, _T_89357}; // @[LoadQueue.scala 191:60:@35841.4]
  assign _T_89359 = conflictPReg_8_5 ? 3'h5 : _T_89358; // @[LoadQueue.scala 191:60:@35842.4]
  assign _T_89360 = conflictPReg_8_6 ? 3'h6 : _T_89359; // @[LoadQueue.scala 191:60:@35843.4]
  assign _T_89361 = conflictPReg_8_7 ? 3'h7 : _T_89360; // @[LoadQueue.scala 191:60:@35844.4]
  assign _T_89362 = conflictPReg_8_8 ? 4'h8 : {{1'd0}, _T_89361}; // @[LoadQueue.scala 191:60:@35845.4]
  assign _T_89363 = conflictPReg_8_9 ? 4'h9 : _T_89362; // @[LoadQueue.scala 191:60:@35846.4]
  assign _T_89364 = conflictPReg_8_10 ? 4'ha : _T_89363; // @[LoadQueue.scala 191:60:@35847.4]
  assign _T_89365 = conflictPReg_8_11 ? 4'hb : _T_89364; // @[LoadQueue.scala 191:60:@35848.4]
  assign _T_89366 = conflictPReg_8_12 ? 4'hc : _T_89365; // @[LoadQueue.scala 191:60:@35849.4]
  assign _T_89367 = conflictPReg_8_13 ? 4'hd : _T_89366; // @[LoadQueue.scala 191:60:@35850.4]
  assign _T_89368 = conflictPReg_8_14 ? 4'he : _T_89367; // @[LoadQueue.scala 191:60:@35851.4]
  assign _T_89369 = conflictPReg_8_15 ? 4'hf : _T_89368; // @[LoadQueue.scala 191:60:@35852.4]
  assign _T_89372 = conflictPReg_8_0 | conflictPReg_8_1; // @[LoadQueue.scala 192:43:@35854.4]
  assign _T_89373 = _T_89372 | conflictPReg_8_2; // @[LoadQueue.scala 192:43:@35855.4]
  assign _T_89374 = _T_89373 | conflictPReg_8_3; // @[LoadQueue.scala 192:43:@35856.4]
  assign _T_89375 = _T_89374 | conflictPReg_8_4; // @[LoadQueue.scala 192:43:@35857.4]
  assign _T_89376 = _T_89375 | conflictPReg_8_5; // @[LoadQueue.scala 192:43:@35858.4]
  assign _T_89377 = _T_89376 | conflictPReg_8_6; // @[LoadQueue.scala 192:43:@35859.4]
  assign _T_89378 = _T_89377 | conflictPReg_8_7; // @[LoadQueue.scala 192:43:@35860.4]
  assign _T_89379 = _T_89378 | conflictPReg_8_8; // @[LoadQueue.scala 192:43:@35861.4]
  assign _T_89380 = _T_89379 | conflictPReg_8_9; // @[LoadQueue.scala 192:43:@35862.4]
  assign _T_89381 = _T_89380 | conflictPReg_8_10; // @[LoadQueue.scala 192:43:@35863.4]
  assign _T_89382 = _T_89381 | conflictPReg_8_11; // @[LoadQueue.scala 192:43:@35864.4]
  assign _T_89383 = _T_89382 | conflictPReg_8_12; // @[LoadQueue.scala 192:43:@35865.4]
  assign _T_89384 = _T_89383 | conflictPReg_8_13; // @[LoadQueue.scala 192:43:@35866.4]
  assign _T_89385 = _T_89384 | conflictPReg_8_14; // @[LoadQueue.scala 192:43:@35867.4]
  assign _T_89386 = _T_89385 | conflictPReg_8_15; // @[LoadQueue.scala 192:43:@35868.4]
  assign _GEN_1392 = 4'h0 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1393 = 4'h1 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1394 = 4'h2 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1395 = 4'h3 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1396 = 4'h4 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1397 = 4'h5 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1398 = 4'h6 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1399 = 4'h7 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1400 = 4'h8 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1401 = 4'h9 == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1402 = 4'ha == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1403 = 4'hb == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1404 = 4'hc == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1405 = 4'hd == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1406 = 4'he == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1407 = 4'hf == _T_89369; // @[LoadQueue.scala 193:43:@35870.6]
  assign _GEN_1409 = 4'h1 == _T_89369 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1410 = 4'h2 == _T_89369 ? shiftedStoreDataKnownPReg_2 : _GEN_1409; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1411 = 4'h3 == _T_89369 ? shiftedStoreDataKnownPReg_3 : _GEN_1410; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1412 = 4'h4 == _T_89369 ? shiftedStoreDataKnownPReg_4 : _GEN_1411; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1413 = 4'h5 == _T_89369 ? shiftedStoreDataKnownPReg_5 : _GEN_1412; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1414 = 4'h6 == _T_89369 ? shiftedStoreDataKnownPReg_6 : _GEN_1413; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1415 = 4'h7 == _T_89369 ? shiftedStoreDataKnownPReg_7 : _GEN_1414; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1416 = 4'h8 == _T_89369 ? shiftedStoreDataKnownPReg_8 : _GEN_1415; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1417 = 4'h9 == _T_89369 ? shiftedStoreDataKnownPReg_9 : _GEN_1416; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1418 = 4'ha == _T_89369 ? shiftedStoreDataKnownPReg_10 : _GEN_1417; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1419 = 4'hb == _T_89369 ? shiftedStoreDataKnownPReg_11 : _GEN_1418; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1420 = 4'hc == _T_89369 ? shiftedStoreDataKnownPReg_12 : _GEN_1419; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1421 = 4'hd == _T_89369 ? shiftedStoreDataKnownPReg_13 : _GEN_1420; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1422 = 4'he == _T_89369 ? shiftedStoreDataKnownPReg_14 : _GEN_1421; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1423 = 4'hf == _T_89369 ? shiftedStoreDataKnownPReg_15 : _GEN_1422; // @[LoadQueue.scala 194:31:@35871.6]
  assign _GEN_1425 = 4'h1 == _T_89369 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1426 = 4'h2 == _T_89369 ? shiftedStoreDataQPreg_2 : _GEN_1425; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1427 = 4'h3 == _T_89369 ? shiftedStoreDataQPreg_3 : _GEN_1426; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1428 = 4'h4 == _T_89369 ? shiftedStoreDataQPreg_4 : _GEN_1427; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1429 = 4'h5 == _T_89369 ? shiftedStoreDataQPreg_5 : _GEN_1428; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1430 = 4'h6 == _T_89369 ? shiftedStoreDataQPreg_6 : _GEN_1429; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1431 = 4'h7 == _T_89369 ? shiftedStoreDataQPreg_7 : _GEN_1430; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1432 = 4'h8 == _T_89369 ? shiftedStoreDataQPreg_8 : _GEN_1431; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1433 = 4'h9 == _T_89369 ? shiftedStoreDataQPreg_9 : _GEN_1432; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1434 = 4'ha == _T_89369 ? shiftedStoreDataQPreg_10 : _GEN_1433; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1435 = 4'hb == _T_89369 ? shiftedStoreDataQPreg_11 : _GEN_1434; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1436 = 4'hc == _T_89369 ? shiftedStoreDataQPreg_12 : _GEN_1435; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1437 = 4'hd == _T_89369 ? shiftedStoreDataQPreg_13 : _GEN_1436; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1438 = 4'he == _T_89369 ? shiftedStoreDataQPreg_14 : _GEN_1437; // @[LoadQueue.scala 195:31:@35872.6]
  assign _GEN_1439 = 4'hf == _T_89369 ? shiftedStoreDataQPreg_15 : _GEN_1438; // @[LoadQueue.scala 195:31:@35872.6]
  assign lastConflict_8_0 = _T_89386 ? _GEN_1392 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_1 = _T_89386 ? _GEN_1393 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_2 = _T_89386 ? _GEN_1394 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_3 = _T_89386 ? _GEN_1395 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_4 = _T_89386 ? _GEN_1396 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_5 = _T_89386 ? _GEN_1397 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_6 = _T_89386 ? _GEN_1398 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_7 = _T_89386 ? _GEN_1399 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_8 = _T_89386 ? _GEN_1400 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_9 = _T_89386 ? _GEN_1401 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_10 = _T_89386 ? _GEN_1402 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_11 = _T_89386 ? _GEN_1403 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_12 = _T_89386 ? _GEN_1404 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_13 = _T_89386 ? _GEN_1405 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_14 = _T_89386 ? _GEN_1406 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign lastConflict_8_15 = _T_89386 ? _GEN_1407 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign canBypass_8 = _T_89386 ? _GEN_1423 : 1'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign bypassVal_8 = _T_89386 ? _GEN_1439 : 32'h0; // @[LoadQueue.scala 192:53:@35869.4]
  assign _T_89492 = conflictPReg_9_2 ? 2'h2 : {{1'd0}, conflictPReg_9_1}; // @[LoadQueue.scala 191:60:@35926.4]
  assign _T_89493 = conflictPReg_9_3 ? 2'h3 : _T_89492; // @[LoadQueue.scala 191:60:@35927.4]
  assign _T_89494 = conflictPReg_9_4 ? 3'h4 : {{1'd0}, _T_89493}; // @[LoadQueue.scala 191:60:@35928.4]
  assign _T_89495 = conflictPReg_9_5 ? 3'h5 : _T_89494; // @[LoadQueue.scala 191:60:@35929.4]
  assign _T_89496 = conflictPReg_9_6 ? 3'h6 : _T_89495; // @[LoadQueue.scala 191:60:@35930.4]
  assign _T_89497 = conflictPReg_9_7 ? 3'h7 : _T_89496; // @[LoadQueue.scala 191:60:@35931.4]
  assign _T_89498 = conflictPReg_9_8 ? 4'h8 : {{1'd0}, _T_89497}; // @[LoadQueue.scala 191:60:@35932.4]
  assign _T_89499 = conflictPReg_9_9 ? 4'h9 : _T_89498; // @[LoadQueue.scala 191:60:@35933.4]
  assign _T_89500 = conflictPReg_9_10 ? 4'ha : _T_89499; // @[LoadQueue.scala 191:60:@35934.4]
  assign _T_89501 = conflictPReg_9_11 ? 4'hb : _T_89500; // @[LoadQueue.scala 191:60:@35935.4]
  assign _T_89502 = conflictPReg_9_12 ? 4'hc : _T_89501; // @[LoadQueue.scala 191:60:@35936.4]
  assign _T_89503 = conflictPReg_9_13 ? 4'hd : _T_89502; // @[LoadQueue.scala 191:60:@35937.4]
  assign _T_89504 = conflictPReg_9_14 ? 4'he : _T_89503; // @[LoadQueue.scala 191:60:@35938.4]
  assign _T_89505 = conflictPReg_9_15 ? 4'hf : _T_89504; // @[LoadQueue.scala 191:60:@35939.4]
  assign _T_89508 = conflictPReg_9_0 | conflictPReg_9_1; // @[LoadQueue.scala 192:43:@35941.4]
  assign _T_89509 = _T_89508 | conflictPReg_9_2; // @[LoadQueue.scala 192:43:@35942.4]
  assign _T_89510 = _T_89509 | conflictPReg_9_3; // @[LoadQueue.scala 192:43:@35943.4]
  assign _T_89511 = _T_89510 | conflictPReg_9_4; // @[LoadQueue.scala 192:43:@35944.4]
  assign _T_89512 = _T_89511 | conflictPReg_9_5; // @[LoadQueue.scala 192:43:@35945.4]
  assign _T_89513 = _T_89512 | conflictPReg_9_6; // @[LoadQueue.scala 192:43:@35946.4]
  assign _T_89514 = _T_89513 | conflictPReg_9_7; // @[LoadQueue.scala 192:43:@35947.4]
  assign _T_89515 = _T_89514 | conflictPReg_9_8; // @[LoadQueue.scala 192:43:@35948.4]
  assign _T_89516 = _T_89515 | conflictPReg_9_9; // @[LoadQueue.scala 192:43:@35949.4]
  assign _T_89517 = _T_89516 | conflictPReg_9_10; // @[LoadQueue.scala 192:43:@35950.4]
  assign _T_89518 = _T_89517 | conflictPReg_9_11; // @[LoadQueue.scala 192:43:@35951.4]
  assign _T_89519 = _T_89518 | conflictPReg_9_12; // @[LoadQueue.scala 192:43:@35952.4]
  assign _T_89520 = _T_89519 | conflictPReg_9_13; // @[LoadQueue.scala 192:43:@35953.4]
  assign _T_89521 = _T_89520 | conflictPReg_9_14; // @[LoadQueue.scala 192:43:@35954.4]
  assign _T_89522 = _T_89521 | conflictPReg_9_15; // @[LoadQueue.scala 192:43:@35955.4]
  assign _GEN_1458 = 4'h0 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1459 = 4'h1 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1460 = 4'h2 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1461 = 4'h3 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1462 = 4'h4 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1463 = 4'h5 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1464 = 4'h6 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1465 = 4'h7 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1466 = 4'h8 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1467 = 4'h9 == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1468 = 4'ha == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1469 = 4'hb == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1470 = 4'hc == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1471 = 4'hd == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1472 = 4'he == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1473 = 4'hf == _T_89505; // @[LoadQueue.scala 193:43:@35957.6]
  assign _GEN_1475 = 4'h1 == _T_89505 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1476 = 4'h2 == _T_89505 ? shiftedStoreDataKnownPReg_2 : _GEN_1475; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1477 = 4'h3 == _T_89505 ? shiftedStoreDataKnownPReg_3 : _GEN_1476; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1478 = 4'h4 == _T_89505 ? shiftedStoreDataKnownPReg_4 : _GEN_1477; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1479 = 4'h5 == _T_89505 ? shiftedStoreDataKnownPReg_5 : _GEN_1478; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1480 = 4'h6 == _T_89505 ? shiftedStoreDataKnownPReg_6 : _GEN_1479; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1481 = 4'h7 == _T_89505 ? shiftedStoreDataKnownPReg_7 : _GEN_1480; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1482 = 4'h8 == _T_89505 ? shiftedStoreDataKnownPReg_8 : _GEN_1481; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1483 = 4'h9 == _T_89505 ? shiftedStoreDataKnownPReg_9 : _GEN_1482; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1484 = 4'ha == _T_89505 ? shiftedStoreDataKnownPReg_10 : _GEN_1483; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1485 = 4'hb == _T_89505 ? shiftedStoreDataKnownPReg_11 : _GEN_1484; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1486 = 4'hc == _T_89505 ? shiftedStoreDataKnownPReg_12 : _GEN_1485; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1487 = 4'hd == _T_89505 ? shiftedStoreDataKnownPReg_13 : _GEN_1486; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1488 = 4'he == _T_89505 ? shiftedStoreDataKnownPReg_14 : _GEN_1487; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1489 = 4'hf == _T_89505 ? shiftedStoreDataKnownPReg_15 : _GEN_1488; // @[LoadQueue.scala 194:31:@35958.6]
  assign _GEN_1491 = 4'h1 == _T_89505 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1492 = 4'h2 == _T_89505 ? shiftedStoreDataQPreg_2 : _GEN_1491; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1493 = 4'h3 == _T_89505 ? shiftedStoreDataQPreg_3 : _GEN_1492; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1494 = 4'h4 == _T_89505 ? shiftedStoreDataQPreg_4 : _GEN_1493; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1495 = 4'h5 == _T_89505 ? shiftedStoreDataQPreg_5 : _GEN_1494; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1496 = 4'h6 == _T_89505 ? shiftedStoreDataQPreg_6 : _GEN_1495; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1497 = 4'h7 == _T_89505 ? shiftedStoreDataQPreg_7 : _GEN_1496; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1498 = 4'h8 == _T_89505 ? shiftedStoreDataQPreg_8 : _GEN_1497; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1499 = 4'h9 == _T_89505 ? shiftedStoreDataQPreg_9 : _GEN_1498; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1500 = 4'ha == _T_89505 ? shiftedStoreDataQPreg_10 : _GEN_1499; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1501 = 4'hb == _T_89505 ? shiftedStoreDataQPreg_11 : _GEN_1500; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1502 = 4'hc == _T_89505 ? shiftedStoreDataQPreg_12 : _GEN_1501; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1503 = 4'hd == _T_89505 ? shiftedStoreDataQPreg_13 : _GEN_1502; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1504 = 4'he == _T_89505 ? shiftedStoreDataQPreg_14 : _GEN_1503; // @[LoadQueue.scala 195:31:@35959.6]
  assign _GEN_1505 = 4'hf == _T_89505 ? shiftedStoreDataQPreg_15 : _GEN_1504; // @[LoadQueue.scala 195:31:@35959.6]
  assign lastConflict_9_0 = _T_89522 ? _GEN_1458 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_1 = _T_89522 ? _GEN_1459 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_2 = _T_89522 ? _GEN_1460 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_3 = _T_89522 ? _GEN_1461 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_4 = _T_89522 ? _GEN_1462 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_5 = _T_89522 ? _GEN_1463 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_6 = _T_89522 ? _GEN_1464 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_7 = _T_89522 ? _GEN_1465 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_8 = _T_89522 ? _GEN_1466 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_9 = _T_89522 ? _GEN_1467 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_10 = _T_89522 ? _GEN_1468 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_11 = _T_89522 ? _GEN_1469 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_12 = _T_89522 ? _GEN_1470 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_13 = _T_89522 ? _GEN_1471 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_14 = _T_89522 ? _GEN_1472 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign lastConflict_9_15 = _T_89522 ? _GEN_1473 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign canBypass_9 = _T_89522 ? _GEN_1489 : 1'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign bypassVal_9 = _T_89522 ? _GEN_1505 : 32'h0; // @[LoadQueue.scala 192:53:@35956.4]
  assign _T_89628 = conflictPReg_10_2 ? 2'h2 : {{1'd0}, conflictPReg_10_1}; // @[LoadQueue.scala 191:60:@36013.4]
  assign _T_89629 = conflictPReg_10_3 ? 2'h3 : _T_89628; // @[LoadQueue.scala 191:60:@36014.4]
  assign _T_89630 = conflictPReg_10_4 ? 3'h4 : {{1'd0}, _T_89629}; // @[LoadQueue.scala 191:60:@36015.4]
  assign _T_89631 = conflictPReg_10_5 ? 3'h5 : _T_89630; // @[LoadQueue.scala 191:60:@36016.4]
  assign _T_89632 = conflictPReg_10_6 ? 3'h6 : _T_89631; // @[LoadQueue.scala 191:60:@36017.4]
  assign _T_89633 = conflictPReg_10_7 ? 3'h7 : _T_89632; // @[LoadQueue.scala 191:60:@36018.4]
  assign _T_89634 = conflictPReg_10_8 ? 4'h8 : {{1'd0}, _T_89633}; // @[LoadQueue.scala 191:60:@36019.4]
  assign _T_89635 = conflictPReg_10_9 ? 4'h9 : _T_89634; // @[LoadQueue.scala 191:60:@36020.4]
  assign _T_89636 = conflictPReg_10_10 ? 4'ha : _T_89635; // @[LoadQueue.scala 191:60:@36021.4]
  assign _T_89637 = conflictPReg_10_11 ? 4'hb : _T_89636; // @[LoadQueue.scala 191:60:@36022.4]
  assign _T_89638 = conflictPReg_10_12 ? 4'hc : _T_89637; // @[LoadQueue.scala 191:60:@36023.4]
  assign _T_89639 = conflictPReg_10_13 ? 4'hd : _T_89638; // @[LoadQueue.scala 191:60:@36024.4]
  assign _T_89640 = conflictPReg_10_14 ? 4'he : _T_89639; // @[LoadQueue.scala 191:60:@36025.4]
  assign _T_89641 = conflictPReg_10_15 ? 4'hf : _T_89640; // @[LoadQueue.scala 191:60:@36026.4]
  assign _T_89644 = conflictPReg_10_0 | conflictPReg_10_1; // @[LoadQueue.scala 192:43:@36028.4]
  assign _T_89645 = _T_89644 | conflictPReg_10_2; // @[LoadQueue.scala 192:43:@36029.4]
  assign _T_89646 = _T_89645 | conflictPReg_10_3; // @[LoadQueue.scala 192:43:@36030.4]
  assign _T_89647 = _T_89646 | conflictPReg_10_4; // @[LoadQueue.scala 192:43:@36031.4]
  assign _T_89648 = _T_89647 | conflictPReg_10_5; // @[LoadQueue.scala 192:43:@36032.4]
  assign _T_89649 = _T_89648 | conflictPReg_10_6; // @[LoadQueue.scala 192:43:@36033.4]
  assign _T_89650 = _T_89649 | conflictPReg_10_7; // @[LoadQueue.scala 192:43:@36034.4]
  assign _T_89651 = _T_89650 | conflictPReg_10_8; // @[LoadQueue.scala 192:43:@36035.4]
  assign _T_89652 = _T_89651 | conflictPReg_10_9; // @[LoadQueue.scala 192:43:@36036.4]
  assign _T_89653 = _T_89652 | conflictPReg_10_10; // @[LoadQueue.scala 192:43:@36037.4]
  assign _T_89654 = _T_89653 | conflictPReg_10_11; // @[LoadQueue.scala 192:43:@36038.4]
  assign _T_89655 = _T_89654 | conflictPReg_10_12; // @[LoadQueue.scala 192:43:@36039.4]
  assign _T_89656 = _T_89655 | conflictPReg_10_13; // @[LoadQueue.scala 192:43:@36040.4]
  assign _T_89657 = _T_89656 | conflictPReg_10_14; // @[LoadQueue.scala 192:43:@36041.4]
  assign _T_89658 = _T_89657 | conflictPReg_10_15; // @[LoadQueue.scala 192:43:@36042.4]
  assign _GEN_1524 = 4'h0 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1525 = 4'h1 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1526 = 4'h2 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1527 = 4'h3 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1528 = 4'h4 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1529 = 4'h5 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1530 = 4'h6 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1531 = 4'h7 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1532 = 4'h8 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1533 = 4'h9 == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1534 = 4'ha == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1535 = 4'hb == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1536 = 4'hc == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1537 = 4'hd == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1538 = 4'he == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1539 = 4'hf == _T_89641; // @[LoadQueue.scala 193:43:@36044.6]
  assign _GEN_1541 = 4'h1 == _T_89641 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1542 = 4'h2 == _T_89641 ? shiftedStoreDataKnownPReg_2 : _GEN_1541; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1543 = 4'h3 == _T_89641 ? shiftedStoreDataKnownPReg_3 : _GEN_1542; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1544 = 4'h4 == _T_89641 ? shiftedStoreDataKnownPReg_4 : _GEN_1543; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1545 = 4'h5 == _T_89641 ? shiftedStoreDataKnownPReg_5 : _GEN_1544; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1546 = 4'h6 == _T_89641 ? shiftedStoreDataKnownPReg_6 : _GEN_1545; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1547 = 4'h7 == _T_89641 ? shiftedStoreDataKnownPReg_7 : _GEN_1546; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1548 = 4'h8 == _T_89641 ? shiftedStoreDataKnownPReg_8 : _GEN_1547; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1549 = 4'h9 == _T_89641 ? shiftedStoreDataKnownPReg_9 : _GEN_1548; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1550 = 4'ha == _T_89641 ? shiftedStoreDataKnownPReg_10 : _GEN_1549; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1551 = 4'hb == _T_89641 ? shiftedStoreDataKnownPReg_11 : _GEN_1550; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1552 = 4'hc == _T_89641 ? shiftedStoreDataKnownPReg_12 : _GEN_1551; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1553 = 4'hd == _T_89641 ? shiftedStoreDataKnownPReg_13 : _GEN_1552; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1554 = 4'he == _T_89641 ? shiftedStoreDataKnownPReg_14 : _GEN_1553; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1555 = 4'hf == _T_89641 ? shiftedStoreDataKnownPReg_15 : _GEN_1554; // @[LoadQueue.scala 194:31:@36045.6]
  assign _GEN_1557 = 4'h1 == _T_89641 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1558 = 4'h2 == _T_89641 ? shiftedStoreDataQPreg_2 : _GEN_1557; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1559 = 4'h3 == _T_89641 ? shiftedStoreDataQPreg_3 : _GEN_1558; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1560 = 4'h4 == _T_89641 ? shiftedStoreDataQPreg_4 : _GEN_1559; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1561 = 4'h5 == _T_89641 ? shiftedStoreDataQPreg_5 : _GEN_1560; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1562 = 4'h6 == _T_89641 ? shiftedStoreDataQPreg_6 : _GEN_1561; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1563 = 4'h7 == _T_89641 ? shiftedStoreDataQPreg_7 : _GEN_1562; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1564 = 4'h8 == _T_89641 ? shiftedStoreDataQPreg_8 : _GEN_1563; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1565 = 4'h9 == _T_89641 ? shiftedStoreDataQPreg_9 : _GEN_1564; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1566 = 4'ha == _T_89641 ? shiftedStoreDataQPreg_10 : _GEN_1565; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1567 = 4'hb == _T_89641 ? shiftedStoreDataQPreg_11 : _GEN_1566; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1568 = 4'hc == _T_89641 ? shiftedStoreDataQPreg_12 : _GEN_1567; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1569 = 4'hd == _T_89641 ? shiftedStoreDataQPreg_13 : _GEN_1568; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1570 = 4'he == _T_89641 ? shiftedStoreDataQPreg_14 : _GEN_1569; // @[LoadQueue.scala 195:31:@36046.6]
  assign _GEN_1571 = 4'hf == _T_89641 ? shiftedStoreDataQPreg_15 : _GEN_1570; // @[LoadQueue.scala 195:31:@36046.6]
  assign lastConflict_10_0 = _T_89658 ? _GEN_1524 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_1 = _T_89658 ? _GEN_1525 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_2 = _T_89658 ? _GEN_1526 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_3 = _T_89658 ? _GEN_1527 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_4 = _T_89658 ? _GEN_1528 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_5 = _T_89658 ? _GEN_1529 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_6 = _T_89658 ? _GEN_1530 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_7 = _T_89658 ? _GEN_1531 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_8 = _T_89658 ? _GEN_1532 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_9 = _T_89658 ? _GEN_1533 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_10 = _T_89658 ? _GEN_1534 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_11 = _T_89658 ? _GEN_1535 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_12 = _T_89658 ? _GEN_1536 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_13 = _T_89658 ? _GEN_1537 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_14 = _T_89658 ? _GEN_1538 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign lastConflict_10_15 = _T_89658 ? _GEN_1539 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign canBypass_10 = _T_89658 ? _GEN_1555 : 1'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign bypassVal_10 = _T_89658 ? _GEN_1571 : 32'h0; // @[LoadQueue.scala 192:53:@36043.4]
  assign _T_89764 = conflictPReg_11_2 ? 2'h2 : {{1'd0}, conflictPReg_11_1}; // @[LoadQueue.scala 191:60:@36100.4]
  assign _T_89765 = conflictPReg_11_3 ? 2'h3 : _T_89764; // @[LoadQueue.scala 191:60:@36101.4]
  assign _T_89766 = conflictPReg_11_4 ? 3'h4 : {{1'd0}, _T_89765}; // @[LoadQueue.scala 191:60:@36102.4]
  assign _T_89767 = conflictPReg_11_5 ? 3'h5 : _T_89766; // @[LoadQueue.scala 191:60:@36103.4]
  assign _T_89768 = conflictPReg_11_6 ? 3'h6 : _T_89767; // @[LoadQueue.scala 191:60:@36104.4]
  assign _T_89769 = conflictPReg_11_7 ? 3'h7 : _T_89768; // @[LoadQueue.scala 191:60:@36105.4]
  assign _T_89770 = conflictPReg_11_8 ? 4'h8 : {{1'd0}, _T_89769}; // @[LoadQueue.scala 191:60:@36106.4]
  assign _T_89771 = conflictPReg_11_9 ? 4'h9 : _T_89770; // @[LoadQueue.scala 191:60:@36107.4]
  assign _T_89772 = conflictPReg_11_10 ? 4'ha : _T_89771; // @[LoadQueue.scala 191:60:@36108.4]
  assign _T_89773 = conflictPReg_11_11 ? 4'hb : _T_89772; // @[LoadQueue.scala 191:60:@36109.4]
  assign _T_89774 = conflictPReg_11_12 ? 4'hc : _T_89773; // @[LoadQueue.scala 191:60:@36110.4]
  assign _T_89775 = conflictPReg_11_13 ? 4'hd : _T_89774; // @[LoadQueue.scala 191:60:@36111.4]
  assign _T_89776 = conflictPReg_11_14 ? 4'he : _T_89775; // @[LoadQueue.scala 191:60:@36112.4]
  assign _T_89777 = conflictPReg_11_15 ? 4'hf : _T_89776; // @[LoadQueue.scala 191:60:@36113.4]
  assign _T_89780 = conflictPReg_11_0 | conflictPReg_11_1; // @[LoadQueue.scala 192:43:@36115.4]
  assign _T_89781 = _T_89780 | conflictPReg_11_2; // @[LoadQueue.scala 192:43:@36116.4]
  assign _T_89782 = _T_89781 | conflictPReg_11_3; // @[LoadQueue.scala 192:43:@36117.4]
  assign _T_89783 = _T_89782 | conflictPReg_11_4; // @[LoadQueue.scala 192:43:@36118.4]
  assign _T_89784 = _T_89783 | conflictPReg_11_5; // @[LoadQueue.scala 192:43:@36119.4]
  assign _T_89785 = _T_89784 | conflictPReg_11_6; // @[LoadQueue.scala 192:43:@36120.4]
  assign _T_89786 = _T_89785 | conflictPReg_11_7; // @[LoadQueue.scala 192:43:@36121.4]
  assign _T_89787 = _T_89786 | conflictPReg_11_8; // @[LoadQueue.scala 192:43:@36122.4]
  assign _T_89788 = _T_89787 | conflictPReg_11_9; // @[LoadQueue.scala 192:43:@36123.4]
  assign _T_89789 = _T_89788 | conflictPReg_11_10; // @[LoadQueue.scala 192:43:@36124.4]
  assign _T_89790 = _T_89789 | conflictPReg_11_11; // @[LoadQueue.scala 192:43:@36125.4]
  assign _T_89791 = _T_89790 | conflictPReg_11_12; // @[LoadQueue.scala 192:43:@36126.4]
  assign _T_89792 = _T_89791 | conflictPReg_11_13; // @[LoadQueue.scala 192:43:@36127.4]
  assign _T_89793 = _T_89792 | conflictPReg_11_14; // @[LoadQueue.scala 192:43:@36128.4]
  assign _T_89794 = _T_89793 | conflictPReg_11_15; // @[LoadQueue.scala 192:43:@36129.4]
  assign _GEN_1590 = 4'h0 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1591 = 4'h1 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1592 = 4'h2 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1593 = 4'h3 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1594 = 4'h4 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1595 = 4'h5 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1596 = 4'h6 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1597 = 4'h7 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1598 = 4'h8 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1599 = 4'h9 == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1600 = 4'ha == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1601 = 4'hb == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1602 = 4'hc == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1603 = 4'hd == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1604 = 4'he == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1605 = 4'hf == _T_89777; // @[LoadQueue.scala 193:43:@36131.6]
  assign _GEN_1607 = 4'h1 == _T_89777 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1608 = 4'h2 == _T_89777 ? shiftedStoreDataKnownPReg_2 : _GEN_1607; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1609 = 4'h3 == _T_89777 ? shiftedStoreDataKnownPReg_3 : _GEN_1608; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1610 = 4'h4 == _T_89777 ? shiftedStoreDataKnownPReg_4 : _GEN_1609; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1611 = 4'h5 == _T_89777 ? shiftedStoreDataKnownPReg_5 : _GEN_1610; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1612 = 4'h6 == _T_89777 ? shiftedStoreDataKnownPReg_6 : _GEN_1611; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1613 = 4'h7 == _T_89777 ? shiftedStoreDataKnownPReg_7 : _GEN_1612; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1614 = 4'h8 == _T_89777 ? shiftedStoreDataKnownPReg_8 : _GEN_1613; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1615 = 4'h9 == _T_89777 ? shiftedStoreDataKnownPReg_9 : _GEN_1614; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1616 = 4'ha == _T_89777 ? shiftedStoreDataKnownPReg_10 : _GEN_1615; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1617 = 4'hb == _T_89777 ? shiftedStoreDataKnownPReg_11 : _GEN_1616; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1618 = 4'hc == _T_89777 ? shiftedStoreDataKnownPReg_12 : _GEN_1617; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1619 = 4'hd == _T_89777 ? shiftedStoreDataKnownPReg_13 : _GEN_1618; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1620 = 4'he == _T_89777 ? shiftedStoreDataKnownPReg_14 : _GEN_1619; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1621 = 4'hf == _T_89777 ? shiftedStoreDataKnownPReg_15 : _GEN_1620; // @[LoadQueue.scala 194:31:@36132.6]
  assign _GEN_1623 = 4'h1 == _T_89777 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1624 = 4'h2 == _T_89777 ? shiftedStoreDataQPreg_2 : _GEN_1623; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1625 = 4'h3 == _T_89777 ? shiftedStoreDataQPreg_3 : _GEN_1624; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1626 = 4'h4 == _T_89777 ? shiftedStoreDataQPreg_4 : _GEN_1625; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1627 = 4'h5 == _T_89777 ? shiftedStoreDataQPreg_5 : _GEN_1626; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1628 = 4'h6 == _T_89777 ? shiftedStoreDataQPreg_6 : _GEN_1627; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1629 = 4'h7 == _T_89777 ? shiftedStoreDataQPreg_7 : _GEN_1628; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1630 = 4'h8 == _T_89777 ? shiftedStoreDataQPreg_8 : _GEN_1629; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1631 = 4'h9 == _T_89777 ? shiftedStoreDataQPreg_9 : _GEN_1630; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1632 = 4'ha == _T_89777 ? shiftedStoreDataQPreg_10 : _GEN_1631; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1633 = 4'hb == _T_89777 ? shiftedStoreDataQPreg_11 : _GEN_1632; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1634 = 4'hc == _T_89777 ? shiftedStoreDataQPreg_12 : _GEN_1633; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1635 = 4'hd == _T_89777 ? shiftedStoreDataQPreg_13 : _GEN_1634; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1636 = 4'he == _T_89777 ? shiftedStoreDataQPreg_14 : _GEN_1635; // @[LoadQueue.scala 195:31:@36133.6]
  assign _GEN_1637 = 4'hf == _T_89777 ? shiftedStoreDataQPreg_15 : _GEN_1636; // @[LoadQueue.scala 195:31:@36133.6]
  assign lastConflict_11_0 = _T_89794 ? _GEN_1590 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_1 = _T_89794 ? _GEN_1591 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_2 = _T_89794 ? _GEN_1592 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_3 = _T_89794 ? _GEN_1593 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_4 = _T_89794 ? _GEN_1594 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_5 = _T_89794 ? _GEN_1595 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_6 = _T_89794 ? _GEN_1596 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_7 = _T_89794 ? _GEN_1597 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_8 = _T_89794 ? _GEN_1598 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_9 = _T_89794 ? _GEN_1599 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_10 = _T_89794 ? _GEN_1600 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_11 = _T_89794 ? _GEN_1601 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_12 = _T_89794 ? _GEN_1602 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_13 = _T_89794 ? _GEN_1603 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_14 = _T_89794 ? _GEN_1604 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign lastConflict_11_15 = _T_89794 ? _GEN_1605 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign canBypass_11 = _T_89794 ? _GEN_1621 : 1'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign bypassVal_11 = _T_89794 ? _GEN_1637 : 32'h0; // @[LoadQueue.scala 192:53:@36130.4]
  assign _T_89900 = conflictPReg_12_2 ? 2'h2 : {{1'd0}, conflictPReg_12_1}; // @[LoadQueue.scala 191:60:@36187.4]
  assign _T_89901 = conflictPReg_12_3 ? 2'h3 : _T_89900; // @[LoadQueue.scala 191:60:@36188.4]
  assign _T_89902 = conflictPReg_12_4 ? 3'h4 : {{1'd0}, _T_89901}; // @[LoadQueue.scala 191:60:@36189.4]
  assign _T_89903 = conflictPReg_12_5 ? 3'h5 : _T_89902; // @[LoadQueue.scala 191:60:@36190.4]
  assign _T_89904 = conflictPReg_12_6 ? 3'h6 : _T_89903; // @[LoadQueue.scala 191:60:@36191.4]
  assign _T_89905 = conflictPReg_12_7 ? 3'h7 : _T_89904; // @[LoadQueue.scala 191:60:@36192.4]
  assign _T_89906 = conflictPReg_12_8 ? 4'h8 : {{1'd0}, _T_89905}; // @[LoadQueue.scala 191:60:@36193.4]
  assign _T_89907 = conflictPReg_12_9 ? 4'h9 : _T_89906; // @[LoadQueue.scala 191:60:@36194.4]
  assign _T_89908 = conflictPReg_12_10 ? 4'ha : _T_89907; // @[LoadQueue.scala 191:60:@36195.4]
  assign _T_89909 = conflictPReg_12_11 ? 4'hb : _T_89908; // @[LoadQueue.scala 191:60:@36196.4]
  assign _T_89910 = conflictPReg_12_12 ? 4'hc : _T_89909; // @[LoadQueue.scala 191:60:@36197.4]
  assign _T_89911 = conflictPReg_12_13 ? 4'hd : _T_89910; // @[LoadQueue.scala 191:60:@36198.4]
  assign _T_89912 = conflictPReg_12_14 ? 4'he : _T_89911; // @[LoadQueue.scala 191:60:@36199.4]
  assign _T_89913 = conflictPReg_12_15 ? 4'hf : _T_89912; // @[LoadQueue.scala 191:60:@36200.4]
  assign _T_89916 = conflictPReg_12_0 | conflictPReg_12_1; // @[LoadQueue.scala 192:43:@36202.4]
  assign _T_89917 = _T_89916 | conflictPReg_12_2; // @[LoadQueue.scala 192:43:@36203.4]
  assign _T_89918 = _T_89917 | conflictPReg_12_3; // @[LoadQueue.scala 192:43:@36204.4]
  assign _T_89919 = _T_89918 | conflictPReg_12_4; // @[LoadQueue.scala 192:43:@36205.4]
  assign _T_89920 = _T_89919 | conflictPReg_12_5; // @[LoadQueue.scala 192:43:@36206.4]
  assign _T_89921 = _T_89920 | conflictPReg_12_6; // @[LoadQueue.scala 192:43:@36207.4]
  assign _T_89922 = _T_89921 | conflictPReg_12_7; // @[LoadQueue.scala 192:43:@36208.4]
  assign _T_89923 = _T_89922 | conflictPReg_12_8; // @[LoadQueue.scala 192:43:@36209.4]
  assign _T_89924 = _T_89923 | conflictPReg_12_9; // @[LoadQueue.scala 192:43:@36210.4]
  assign _T_89925 = _T_89924 | conflictPReg_12_10; // @[LoadQueue.scala 192:43:@36211.4]
  assign _T_89926 = _T_89925 | conflictPReg_12_11; // @[LoadQueue.scala 192:43:@36212.4]
  assign _T_89927 = _T_89926 | conflictPReg_12_12; // @[LoadQueue.scala 192:43:@36213.4]
  assign _T_89928 = _T_89927 | conflictPReg_12_13; // @[LoadQueue.scala 192:43:@36214.4]
  assign _T_89929 = _T_89928 | conflictPReg_12_14; // @[LoadQueue.scala 192:43:@36215.4]
  assign _T_89930 = _T_89929 | conflictPReg_12_15; // @[LoadQueue.scala 192:43:@36216.4]
  assign _GEN_1656 = 4'h0 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1657 = 4'h1 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1658 = 4'h2 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1659 = 4'h3 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1660 = 4'h4 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1661 = 4'h5 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1662 = 4'h6 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1663 = 4'h7 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1664 = 4'h8 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1665 = 4'h9 == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1666 = 4'ha == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1667 = 4'hb == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1668 = 4'hc == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1669 = 4'hd == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1670 = 4'he == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1671 = 4'hf == _T_89913; // @[LoadQueue.scala 193:43:@36218.6]
  assign _GEN_1673 = 4'h1 == _T_89913 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1674 = 4'h2 == _T_89913 ? shiftedStoreDataKnownPReg_2 : _GEN_1673; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1675 = 4'h3 == _T_89913 ? shiftedStoreDataKnownPReg_3 : _GEN_1674; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1676 = 4'h4 == _T_89913 ? shiftedStoreDataKnownPReg_4 : _GEN_1675; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1677 = 4'h5 == _T_89913 ? shiftedStoreDataKnownPReg_5 : _GEN_1676; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1678 = 4'h6 == _T_89913 ? shiftedStoreDataKnownPReg_6 : _GEN_1677; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1679 = 4'h7 == _T_89913 ? shiftedStoreDataKnownPReg_7 : _GEN_1678; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1680 = 4'h8 == _T_89913 ? shiftedStoreDataKnownPReg_8 : _GEN_1679; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1681 = 4'h9 == _T_89913 ? shiftedStoreDataKnownPReg_9 : _GEN_1680; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1682 = 4'ha == _T_89913 ? shiftedStoreDataKnownPReg_10 : _GEN_1681; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1683 = 4'hb == _T_89913 ? shiftedStoreDataKnownPReg_11 : _GEN_1682; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1684 = 4'hc == _T_89913 ? shiftedStoreDataKnownPReg_12 : _GEN_1683; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1685 = 4'hd == _T_89913 ? shiftedStoreDataKnownPReg_13 : _GEN_1684; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1686 = 4'he == _T_89913 ? shiftedStoreDataKnownPReg_14 : _GEN_1685; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1687 = 4'hf == _T_89913 ? shiftedStoreDataKnownPReg_15 : _GEN_1686; // @[LoadQueue.scala 194:31:@36219.6]
  assign _GEN_1689 = 4'h1 == _T_89913 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1690 = 4'h2 == _T_89913 ? shiftedStoreDataQPreg_2 : _GEN_1689; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1691 = 4'h3 == _T_89913 ? shiftedStoreDataQPreg_3 : _GEN_1690; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1692 = 4'h4 == _T_89913 ? shiftedStoreDataQPreg_4 : _GEN_1691; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1693 = 4'h5 == _T_89913 ? shiftedStoreDataQPreg_5 : _GEN_1692; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1694 = 4'h6 == _T_89913 ? shiftedStoreDataQPreg_6 : _GEN_1693; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1695 = 4'h7 == _T_89913 ? shiftedStoreDataQPreg_7 : _GEN_1694; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1696 = 4'h8 == _T_89913 ? shiftedStoreDataQPreg_8 : _GEN_1695; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1697 = 4'h9 == _T_89913 ? shiftedStoreDataQPreg_9 : _GEN_1696; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1698 = 4'ha == _T_89913 ? shiftedStoreDataQPreg_10 : _GEN_1697; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1699 = 4'hb == _T_89913 ? shiftedStoreDataQPreg_11 : _GEN_1698; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1700 = 4'hc == _T_89913 ? shiftedStoreDataQPreg_12 : _GEN_1699; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1701 = 4'hd == _T_89913 ? shiftedStoreDataQPreg_13 : _GEN_1700; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1702 = 4'he == _T_89913 ? shiftedStoreDataQPreg_14 : _GEN_1701; // @[LoadQueue.scala 195:31:@36220.6]
  assign _GEN_1703 = 4'hf == _T_89913 ? shiftedStoreDataQPreg_15 : _GEN_1702; // @[LoadQueue.scala 195:31:@36220.6]
  assign lastConflict_12_0 = _T_89930 ? _GEN_1656 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_1 = _T_89930 ? _GEN_1657 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_2 = _T_89930 ? _GEN_1658 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_3 = _T_89930 ? _GEN_1659 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_4 = _T_89930 ? _GEN_1660 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_5 = _T_89930 ? _GEN_1661 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_6 = _T_89930 ? _GEN_1662 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_7 = _T_89930 ? _GEN_1663 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_8 = _T_89930 ? _GEN_1664 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_9 = _T_89930 ? _GEN_1665 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_10 = _T_89930 ? _GEN_1666 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_11 = _T_89930 ? _GEN_1667 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_12 = _T_89930 ? _GEN_1668 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_13 = _T_89930 ? _GEN_1669 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_14 = _T_89930 ? _GEN_1670 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign lastConflict_12_15 = _T_89930 ? _GEN_1671 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign canBypass_12 = _T_89930 ? _GEN_1687 : 1'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign bypassVal_12 = _T_89930 ? _GEN_1703 : 32'h0; // @[LoadQueue.scala 192:53:@36217.4]
  assign _T_90036 = conflictPReg_13_2 ? 2'h2 : {{1'd0}, conflictPReg_13_1}; // @[LoadQueue.scala 191:60:@36274.4]
  assign _T_90037 = conflictPReg_13_3 ? 2'h3 : _T_90036; // @[LoadQueue.scala 191:60:@36275.4]
  assign _T_90038 = conflictPReg_13_4 ? 3'h4 : {{1'd0}, _T_90037}; // @[LoadQueue.scala 191:60:@36276.4]
  assign _T_90039 = conflictPReg_13_5 ? 3'h5 : _T_90038; // @[LoadQueue.scala 191:60:@36277.4]
  assign _T_90040 = conflictPReg_13_6 ? 3'h6 : _T_90039; // @[LoadQueue.scala 191:60:@36278.4]
  assign _T_90041 = conflictPReg_13_7 ? 3'h7 : _T_90040; // @[LoadQueue.scala 191:60:@36279.4]
  assign _T_90042 = conflictPReg_13_8 ? 4'h8 : {{1'd0}, _T_90041}; // @[LoadQueue.scala 191:60:@36280.4]
  assign _T_90043 = conflictPReg_13_9 ? 4'h9 : _T_90042; // @[LoadQueue.scala 191:60:@36281.4]
  assign _T_90044 = conflictPReg_13_10 ? 4'ha : _T_90043; // @[LoadQueue.scala 191:60:@36282.4]
  assign _T_90045 = conflictPReg_13_11 ? 4'hb : _T_90044; // @[LoadQueue.scala 191:60:@36283.4]
  assign _T_90046 = conflictPReg_13_12 ? 4'hc : _T_90045; // @[LoadQueue.scala 191:60:@36284.4]
  assign _T_90047 = conflictPReg_13_13 ? 4'hd : _T_90046; // @[LoadQueue.scala 191:60:@36285.4]
  assign _T_90048 = conflictPReg_13_14 ? 4'he : _T_90047; // @[LoadQueue.scala 191:60:@36286.4]
  assign _T_90049 = conflictPReg_13_15 ? 4'hf : _T_90048; // @[LoadQueue.scala 191:60:@36287.4]
  assign _T_90052 = conflictPReg_13_0 | conflictPReg_13_1; // @[LoadQueue.scala 192:43:@36289.4]
  assign _T_90053 = _T_90052 | conflictPReg_13_2; // @[LoadQueue.scala 192:43:@36290.4]
  assign _T_90054 = _T_90053 | conflictPReg_13_3; // @[LoadQueue.scala 192:43:@36291.4]
  assign _T_90055 = _T_90054 | conflictPReg_13_4; // @[LoadQueue.scala 192:43:@36292.4]
  assign _T_90056 = _T_90055 | conflictPReg_13_5; // @[LoadQueue.scala 192:43:@36293.4]
  assign _T_90057 = _T_90056 | conflictPReg_13_6; // @[LoadQueue.scala 192:43:@36294.4]
  assign _T_90058 = _T_90057 | conflictPReg_13_7; // @[LoadQueue.scala 192:43:@36295.4]
  assign _T_90059 = _T_90058 | conflictPReg_13_8; // @[LoadQueue.scala 192:43:@36296.4]
  assign _T_90060 = _T_90059 | conflictPReg_13_9; // @[LoadQueue.scala 192:43:@36297.4]
  assign _T_90061 = _T_90060 | conflictPReg_13_10; // @[LoadQueue.scala 192:43:@36298.4]
  assign _T_90062 = _T_90061 | conflictPReg_13_11; // @[LoadQueue.scala 192:43:@36299.4]
  assign _T_90063 = _T_90062 | conflictPReg_13_12; // @[LoadQueue.scala 192:43:@36300.4]
  assign _T_90064 = _T_90063 | conflictPReg_13_13; // @[LoadQueue.scala 192:43:@36301.4]
  assign _T_90065 = _T_90064 | conflictPReg_13_14; // @[LoadQueue.scala 192:43:@36302.4]
  assign _T_90066 = _T_90065 | conflictPReg_13_15; // @[LoadQueue.scala 192:43:@36303.4]
  assign _GEN_1722 = 4'h0 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1723 = 4'h1 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1724 = 4'h2 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1725 = 4'h3 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1726 = 4'h4 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1727 = 4'h5 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1728 = 4'h6 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1729 = 4'h7 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1730 = 4'h8 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1731 = 4'h9 == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1732 = 4'ha == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1733 = 4'hb == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1734 = 4'hc == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1735 = 4'hd == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1736 = 4'he == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1737 = 4'hf == _T_90049; // @[LoadQueue.scala 193:43:@36305.6]
  assign _GEN_1739 = 4'h1 == _T_90049 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1740 = 4'h2 == _T_90049 ? shiftedStoreDataKnownPReg_2 : _GEN_1739; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1741 = 4'h3 == _T_90049 ? shiftedStoreDataKnownPReg_3 : _GEN_1740; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1742 = 4'h4 == _T_90049 ? shiftedStoreDataKnownPReg_4 : _GEN_1741; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1743 = 4'h5 == _T_90049 ? shiftedStoreDataKnownPReg_5 : _GEN_1742; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1744 = 4'h6 == _T_90049 ? shiftedStoreDataKnownPReg_6 : _GEN_1743; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1745 = 4'h7 == _T_90049 ? shiftedStoreDataKnownPReg_7 : _GEN_1744; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1746 = 4'h8 == _T_90049 ? shiftedStoreDataKnownPReg_8 : _GEN_1745; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1747 = 4'h9 == _T_90049 ? shiftedStoreDataKnownPReg_9 : _GEN_1746; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1748 = 4'ha == _T_90049 ? shiftedStoreDataKnownPReg_10 : _GEN_1747; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1749 = 4'hb == _T_90049 ? shiftedStoreDataKnownPReg_11 : _GEN_1748; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1750 = 4'hc == _T_90049 ? shiftedStoreDataKnownPReg_12 : _GEN_1749; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1751 = 4'hd == _T_90049 ? shiftedStoreDataKnownPReg_13 : _GEN_1750; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1752 = 4'he == _T_90049 ? shiftedStoreDataKnownPReg_14 : _GEN_1751; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1753 = 4'hf == _T_90049 ? shiftedStoreDataKnownPReg_15 : _GEN_1752; // @[LoadQueue.scala 194:31:@36306.6]
  assign _GEN_1755 = 4'h1 == _T_90049 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1756 = 4'h2 == _T_90049 ? shiftedStoreDataQPreg_2 : _GEN_1755; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1757 = 4'h3 == _T_90049 ? shiftedStoreDataQPreg_3 : _GEN_1756; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1758 = 4'h4 == _T_90049 ? shiftedStoreDataQPreg_4 : _GEN_1757; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1759 = 4'h5 == _T_90049 ? shiftedStoreDataQPreg_5 : _GEN_1758; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1760 = 4'h6 == _T_90049 ? shiftedStoreDataQPreg_6 : _GEN_1759; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1761 = 4'h7 == _T_90049 ? shiftedStoreDataQPreg_7 : _GEN_1760; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1762 = 4'h8 == _T_90049 ? shiftedStoreDataQPreg_8 : _GEN_1761; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1763 = 4'h9 == _T_90049 ? shiftedStoreDataQPreg_9 : _GEN_1762; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1764 = 4'ha == _T_90049 ? shiftedStoreDataQPreg_10 : _GEN_1763; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1765 = 4'hb == _T_90049 ? shiftedStoreDataQPreg_11 : _GEN_1764; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1766 = 4'hc == _T_90049 ? shiftedStoreDataQPreg_12 : _GEN_1765; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1767 = 4'hd == _T_90049 ? shiftedStoreDataQPreg_13 : _GEN_1766; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1768 = 4'he == _T_90049 ? shiftedStoreDataQPreg_14 : _GEN_1767; // @[LoadQueue.scala 195:31:@36307.6]
  assign _GEN_1769 = 4'hf == _T_90049 ? shiftedStoreDataQPreg_15 : _GEN_1768; // @[LoadQueue.scala 195:31:@36307.6]
  assign lastConflict_13_0 = _T_90066 ? _GEN_1722 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_1 = _T_90066 ? _GEN_1723 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_2 = _T_90066 ? _GEN_1724 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_3 = _T_90066 ? _GEN_1725 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_4 = _T_90066 ? _GEN_1726 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_5 = _T_90066 ? _GEN_1727 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_6 = _T_90066 ? _GEN_1728 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_7 = _T_90066 ? _GEN_1729 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_8 = _T_90066 ? _GEN_1730 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_9 = _T_90066 ? _GEN_1731 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_10 = _T_90066 ? _GEN_1732 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_11 = _T_90066 ? _GEN_1733 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_12 = _T_90066 ? _GEN_1734 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_13 = _T_90066 ? _GEN_1735 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_14 = _T_90066 ? _GEN_1736 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign lastConflict_13_15 = _T_90066 ? _GEN_1737 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign canBypass_13 = _T_90066 ? _GEN_1753 : 1'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign bypassVal_13 = _T_90066 ? _GEN_1769 : 32'h0; // @[LoadQueue.scala 192:53:@36304.4]
  assign _T_90172 = conflictPReg_14_2 ? 2'h2 : {{1'd0}, conflictPReg_14_1}; // @[LoadQueue.scala 191:60:@36361.4]
  assign _T_90173 = conflictPReg_14_3 ? 2'h3 : _T_90172; // @[LoadQueue.scala 191:60:@36362.4]
  assign _T_90174 = conflictPReg_14_4 ? 3'h4 : {{1'd0}, _T_90173}; // @[LoadQueue.scala 191:60:@36363.4]
  assign _T_90175 = conflictPReg_14_5 ? 3'h5 : _T_90174; // @[LoadQueue.scala 191:60:@36364.4]
  assign _T_90176 = conflictPReg_14_6 ? 3'h6 : _T_90175; // @[LoadQueue.scala 191:60:@36365.4]
  assign _T_90177 = conflictPReg_14_7 ? 3'h7 : _T_90176; // @[LoadQueue.scala 191:60:@36366.4]
  assign _T_90178 = conflictPReg_14_8 ? 4'h8 : {{1'd0}, _T_90177}; // @[LoadQueue.scala 191:60:@36367.4]
  assign _T_90179 = conflictPReg_14_9 ? 4'h9 : _T_90178; // @[LoadQueue.scala 191:60:@36368.4]
  assign _T_90180 = conflictPReg_14_10 ? 4'ha : _T_90179; // @[LoadQueue.scala 191:60:@36369.4]
  assign _T_90181 = conflictPReg_14_11 ? 4'hb : _T_90180; // @[LoadQueue.scala 191:60:@36370.4]
  assign _T_90182 = conflictPReg_14_12 ? 4'hc : _T_90181; // @[LoadQueue.scala 191:60:@36371.4]
  assign _T_90183 = conflictPReg_14_13 ? 4'hd : _T_90182; // @[LoadQueue.scala 191:60:@36372.4]
  assign _T_90184 = conflictPReg_14_14 ? 4'he : _T_90183; // @[LoadQueue.scala 191:60:@36373.4]
  assign _T_90185 = conflictPReg_14_15 ? 4'hf : _T_90184; // @[LoadQueue.scala 191:60:@36374.4]
  assign _T_90188 = conflictPReg_14_0 | conflictPReg_14_1; // @[LoadQueue.scala 192:43:@36376.4]
  assign _T_90189 = _T_90188 | conflictPReg_14_2; // @[LoadQueue.scala 192:43:@36377.4]
  assign _T_90190 = _T_90189 | conflictPReg_14_3; // @[LoadQueue.scala 192:43:@36378.4]
  assign _T_90191 = _T_90190 | conflictPReg_14_4; // @[LoadQueue.scala 192:43:@36379.4]
  assign _T_90192 = _T_90191 | conflictPReg_14_5; // @[LoadQueue.scala 192:43:@36380.4]
  assign _T_90193 = _T_90192 | conflictPReg_14_6; // @[LoadQueue.scala 192:43:@36381.4]
  assign _T_90194 = _T_90193 | conflictPReg_14_7; // @[LoadQueue.scala 192:43:@36382.4]
  assign _T_90195 = _T_90194 | conflictPReg_14_8; // @[LoadQueue.scala 192:43:@36383.4]
  assign _T_90196 = _T_90195 | conflictPReg_14_9; // @[LoadQueue.scala 192:43:@36384.4]
  assign _T_90197 = _T_90196 | conflictPReg_14_10; // @[LoadQueue.scala 192:43:@36385.4]
  assign _T_90198 = _T_90197 | conflictPReg_14_11; // @[LoadQueue.scala 192:43:@36386.4]
  assign _T_90199 = _T_90198 | conflictPReg_14_12; // @[LoadQueue.scala 192:43:@36387.4]
  assign _T_90200 = _T_90199 | conflictPReg_14_13; // @[LoadQueue.scala 192:43:@36388.4]
  assign _T_90201 = _T_90200 | conflictPReg_14_14; // @[LoadQueue.scala 192:43:@36389.4]
  assign _T_90202 = _T_90201 | conflictPReg_14_15; // @[LoadQueue.scala 192:43:@36390.4]
  assign _GEN_1788 = 4'h0 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1789 = 4'h1 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1790 = 4'h2 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1791 = 4'h3 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1792 = 4'h4 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1793 = 4'h5 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1794 = 4'h6 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1795 = 4'h7 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1796 = 4'h8 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1797 = 4'h9 == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1798 = 4'ha == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1799 = 4'hb == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1800 = 4'hc == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1801 = 4'hd == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1802 = 4'he == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1803 = 4'hf == _T_90185; // @[LoadQueue.scala 193:43:@36392.6]
  assign _GEN_1805 = 4'h1 == _T_90185 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1806 = 4'h2 == _T_90185 ? shiftedStoreDataKnownPReg_2 : _GEN_1805; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1807 = 4'h3 == _T_90185 ? shiftedStoreDataKnownPReg_3 : _GEN_1806; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1808 = 4'h4 == _T_90185 ? shiftedStoreDataKnownPReg_4 : _GEN_1807; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1809 = 4'h5 == _T_90185 ? shiftedStoreDataKnownPReg_5 : _GEN_1808; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1810 = 4'h6 == _T_90185 ? shiftedStoreDataKnownPReg_6 : _GEN_1809; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1811 = 4'h7 == _T_90185 ? shiftedStoreDataKnownPReg_7 : _GEN_1810; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1812 = 4'h8 == _T_90185 ? shiftedStoreDataKnownPReg_8 : _GEN_1811; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1813 = 4'h9 == _T_90185 ? shiftedStoreDataKnownPReg_9 : _GEN_1812; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1814 = 4'ha == _T_90185 ? shiftedStoreDataKnownPReg_10 : _GEN_1813; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1815 = 4'hb == _T_90185 ? shiftedStoreDataKnownPReg_11 : _GEN_1814; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1816 = 4'hc == _T_90185 ? shiftedStoreDataKnownPReg_12 : _GEN_1815; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1817 = 4'hd == _T_90185 ? shiftedStoreDataKnownPReg_13 : _GEN_1816; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1818 = 4'he == _T_90185 ? shiftedStoreDataKnownPReg_14 : _GEN_1817; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1819 = 4'hf == _T_90185 ? shiftedStoreDataKnownPReg_15 : _GEN_1818; // @[LoadQueue.scala 194:31:@36393.6]
  assign _GEN_1821 = 4'h1 == _T_90185 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1822 = 4'h2 == _T_90185 ? shiftedStoreDataQPreg_2 : _GEN_1821; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1823 = 4'h3 == _T_90185 ? shiftedStoreDataQPreg_3 : _GEN_1822; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1824 = 4'h4 == _T_90185 ? shiftedStoreDataQPreg_4 : _GEN_1823; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1825 = 4'h5 == _T_90185 ? shiftedStoreDataQPreg_5 : _GEN_1824; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1826 = 4'h6 == _T_90185 ? shiftedStoreDataQPreg_6 : _GEN_1825; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1827 = 4'h7 == _T_90185 ? shiftedStoreDataQPreg_7 : _GEN_1826; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1828 = 4'h8 == _T_90185 ? shiftedStoreDataQPreg_8 : _GEN_1827; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1829 = 4'h9 == _T_90185 ? shiftedStoreDataQPreg_9 : _GEN_1828; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1830 = 4'ha == _T_90185 ? shiftedStoreDataQPreg_10 : _GEN_1829; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1831 = 4'hb == _T_90185 ? shiftedStoreDataQPreg_11 : _GEN_1830; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1832 = 4'hc == _T_90185 ? shiftedStoreDataQPreg_12 : _GEN_1831; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1833 = 4'hd == _T_90185 ? shiftedStoreDataQPreg_13 : _GEN_1832; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1834 = 4'he == _T_90185 ? shiftedStoreDataQPreg_14 : _GEN_1833; // @[LoadQueue.scala 195:31:@36394.6]
  assign _GEN_1835 = 4'hf == _T_90185 ? shiftedStoreDataQPreg_15 : _GEN_1834; // @[LoadQueue.scala 195:31:@36394.6]
  assign lastConflict_14_0 = _T_90202 ? _GEN_1788 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_1 = _T_90202 ? _GEN_1789 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_2 = _T_90202 ? _GEN_1790 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_3 = _T_90202 ? _GEN_1791 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_4 = _T_90202 ? _GEN_1792 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_5 = _T_90202 ? _GEN_1793 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_6 = _T_90202 ? _GEN_1794 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_7 = _T_90202 ? _GEN_1795 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_8 = _T_90202 ? _GEN_1796 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_9 = _T_90202 ? _GEN_1797 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_10 = _T_90202 ? _GEN_1798 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_11 = _T_90202 ? _GEN_1799 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_12 = _T_90202 ? _GEN_1800 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_13 = _T_90202 ? _GEN_1801 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_14 = _T_90202 ? _GEN_1802 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign lastConflict_14_15 = _T_90202 ? _GEN_1803 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign canBypass_14 = _T_90202 ? _GEN_1819 : 1'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign bypassVal_14 = _T_90202 ? _GEN_1835 : 32'h0; // @[LoadQueue.scala 192:53:@36391.4]
  assign _T_90308 = conflictPReg_15_2 ? 2'h2 : {{1'd0}, conflictPReg_15_1}; // @[LoadQueue.scala 191:60:@36448.4]
  assign _T_90309 = conflictPReg_15_3 ? 2'h3 : _T_90308; // @[LoadQueue.scala 191:60:@36449.4]
  assign _T_90310 = conflictPReg_15_4 ? 3'h4 : {{1'd0}, _T_90309}; // @[LoadQueue.scala 191:60:@36450.4]
  assign _T_90311 = conflictPReg_15_5 ? 3'h5 : _T_90310; // @[LoadQueue.scala 191:60:@36451.4]
  assign _T_90312 = conflictPReg_15_6 ? 3'h6 : _T_90311; // @[LoadQueue.scala 191:60:@36452.4]
  assign _T_90313 = conflictPReg_15_7 ? 3'h7 : _T_90312; // @[LoadQueue.scala 191:60:@36453.4]
  assign _T_90314 = conflictPReg_15_8 ? 4'h8 : {{1'd0}, _T_90313}; // @[LoadQueue.scala 191:60:@36454.4]
  assign _T_90315 = conflictPReg_15_9 ? 4'h9 : _T_90314; // @[LoadQueue.scala 191:60:@36455.4]
  assign _T_90316 = conflictPReg_15_10 ? 4'ha : _T_90315; // @[LoadQueue.scala 191:60:@36456.4]
  assign _T_90317 = conflictPReg_15_11 ? 4'hb : _T_90316; // @[LoadQueue.scala 191:60:@36457.4]
  assign _T_90318 = conflictPReg_15_12 ? 4'hc : _T_90317; // @[LoadQueue.scala 191:60:@36458.4]
  assign _T_90319 = conflictPReg_15_13 ? 4'hd : _T_90318; // @[LoadQueue.scala 191:60:@36459.4]
  assign _T_90320 = conflictPReg_15_14 ? 4'he : _T_90319; // @[LoadQueue.scala 191:60:@36460.4]
  assign _T_90321 = conflictPReg_15_15 ? 4'hf : _T_90320; // @[LoadQueue.scala 191:60:@36461.4]
  assign _T_90324 = conflictPReg_15_0 | conflictPReg_15_1; // @[LoadQueue.scala 192:43:@36463.4]
  assign _T_90325 = _T_90324 | conflictPReg_15_2; // @[LoadQueue.scala 192:43:@36464.4]
  assign _T_90326 = _T_90325 | conflictPReg_15_3; // @[LoadQueue.scala 192:43:@36465.4]
  assign _T_90327 = _T_90326 | conflictPReg_15_4; // @[LoadQueue.scala 192:43:@36466.4]
  assign _T_90328 = _T_90327 | conflictPReg_15_5; // @[LoadQueue.scala 192:43:@36467.4]
  assign _T_90329 = _T_90328 | conflictPReg_15_6; // @[LoadQueue.scala 192:43:@36468.4]
  assign _T_90330 = _T_90329 | conflictPReg_15_7; // @[LoadQueue.scala 192:43:@36469.4]
  assign _T_90331 = _T_90330 | conflictPReg_15_8; // @[LoadQueue.scala 192:43:@36470.4]
  assign _T_90332 = _T_90331 | conflictPReg_15_9; // @[LoadQueue.scala 192:43:@36471.4]
  assign _T_90333 = _T_90332 | conflictPReg_15_10; // @[LoadQueue.scala 192:43:@36472.4]
  assign _T_90334 = _T_90333 | conflictPReg_15_11; // @[LoadQueue.scala 192:43:@36473.4]
  assign _T_90335 = _T_90334 | conflictPReg_15_12; // @[LoadQueue.scala 192:43:@36474.4]
  assign _T_90336 = _T_90335 | conflictPReg_15_13; // @[LoadQueue.scala 192:43:@36475.4]
  assign _T_90337 = _T_90336 | conflictPReg_15_14; // @[LoadQueue.scala 192:43:@36476.4]
  assign _T_90338 = _T_90337 | conflictPReg_15_15; // @[LoadQueue.scala 192:43:@36477.4]
  assign _GEN_1854 = 4'h0 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1855 = 4'h1 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1856 = 4'h2 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1857 = 4'h3 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1858 = 4'h4 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1859 = 4'h5 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1860 = 4'h6 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1861 = 4'h7 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1862 = 4'h8 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1863 = 4'h9 == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1864 = 4'ha == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1865 = 4'hb == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1866 = 4'hc == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1867 = 4'hd == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1868 = 4'he == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1869 = 4'hf == _T_90321; // @[LoadQueue.scala 193:43:@36479.6]
  assign _GEN_1871 = 4'h1 == _T_90321 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1872 = 4'h2 == _T_90321 ? shiftedStoreDataKnownPReg_2 : _GEN_1871; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1873 = 4'h3 == _T_90321 ? shiftedStoreDataKnownPReg_3 : _GEN_1872; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1874 = 4'h4 == _T_90321 ? shiftedStoreDataKnownPReg_4 : _GEN_1873; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1875 = 4'h5 == _T_90321 ? shiftedStoreDataKnownPReg_5 : _GEN_1874; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1876 = 4'h6 == _T_90321 ? shiftedStoreDataKnownPReg_6 : _GEN_1875; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1877 = 4'h7 == _T_90321 ? shiftedStoreDataKnownPReg_7 : _GEN_1876; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1878 = 4'h8 == _T_90321 ? shiftedStoreDataKnownPReg_8 : _GEN_1877; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1879 = 4'h9 == _T_90321 ? shiftedStoreDataKnownPReg_9 : _GEN_1878; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1880 = 4'ha == _T_90321 ? shiftedStoreDataKnownPReg_10 : _GEN_1879; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1881 = 4'hb == _T_90321 ? shiftedStoreDataKnownPReg_11 : _GEN_1880; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1882 = 4'hc == _T_90321 ? shiftedStoreDataKnownPReg_12 : _GEN_1881; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1883 = 4'hd == _T_90321 ? shiftedStoreDataKnownPReg_13 : _GEN_1882; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1884 = 4'he == _T_90321 ? shiftedStoreDataKnownPReg_14 : _GEN_1883; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1885 = 4'hf == _T_90321 ? shiftedStoreDataKnownPReg_15 : _GEN_1884; // @[LoadQueue.scala 194:31:@36480.6]
  assign _GEN_1887 = 4'h1 == _T_90321 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1888 = 4'h2 == _T_90321 ? shiftedStoreDataQPreg_2 : _GEN_1887; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1889 = 4'h3 == _T_90321 ? shiftedStoreDataQPreg_3 : _GEN_1888; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1890 = 4'h4 == _T_90321 ? shiftedStoreDataQPreg_4 : _GEN_1889; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1891 = 4'h5 == _T_90321 ? shiftedStoreDataQPreg_5 : _GEN_1890; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1892 = 4'h6 == _T_90321 ? shiftedStoreDataQPreg_6 : _GEN_1891; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1893 = 4'h7 == _T_90321 ? shiftedStoreDataQPreg_7 : _GEN_1892; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1894 = 4'h8 == _T_90321 ? shiftedStoreDataQPreg_8 : _GEN_1893; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1895 = 4'h9 == _T_90321 ? shiftedStoreDataQPreg_9 : _GEN_1894; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1896 = 4'ha == _T_90321 ? shiftedStoreDataQPreg_10 : _GEN_1895; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1897 = 4'hb == _T_90321 ? shiftedStoreDataQPreg_11 : _GEN_1896; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1898 = 4'hc == _T_90321 ? shiftedStoreDataQPreg_12 : _GEN_1897; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1899 = 4'hd == _T_90321 ? shiftedStoreDataQPreg_13 : _GEN_1898; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1900 = 4'he == _T_90321 ? shiftedStoreDataQPreg_14 : _GEN_1899; // @[LoadQueue.scala 195:31:@36481.6]
  assign _GEN_1901 = 4'hf == _T_90321 ? shiftedStoreDataQPreg_15 : _GEN_1900; // @[LoadQueue.scala 195:31:@36481.6]
  assign lastConflict_15_0 = _T_90338 ? _GEN_1854 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_1 = _T_90338 ? _GEN_1855 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_2 = _T_90338 ? _GEN_1856 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_3 = _T_90338 ? _GEN_1857 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_4 = _T_90338 ? _GEN_1858 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_5 = _T_90338 ? _GEN_1859 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_6 = _T_90338 ? _GEN_1860 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_7 = _T_90338 ? _GEN_1861 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_8 = _T_90338 ? _GEN_1862 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_9 = _T_90338 ? _GEN_1863 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_10 = _T_90338 ? _GEN_1864 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_11 = _T_90338 ? _GEN_1865 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_12 = _T_90338 ? _GEN_1866 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_13 = _T_90338 ? _GEN_1867 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_14 = _T_90338 ? _GEN_1868 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign lastConflict_15_15 = _T_90338 ? _GEN_1869 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign canBypass_15 = _T_90338 ? _GEN_1885 : 1'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign bypassVal_15 = _T_90338 ? _GEN_1901 : 32'h0; // @[LoadQueue.scala 192:53:@36478.4]
  assign _T_90398 = 16'h1 << head; // @[OneHot.scala 52:12:@36486.4]
  assign _T_90400 = _T_90398[0]; // @[util.scala 33:60:@36488.4]
  assign _T_90401 = _T_90398[1]; // @[util.scala 33:60:@36489.4]
  assign _T_90402 = _T_90398[2]; // @[util.scala 33:60:@36490.4]
  assign _T_90403 = _T_90398[3]; // @[util.scala 33:60:@36491.4]
  assign _T_90404 = _T_90398[4]; // @[util.scala 33:60:@36492.4]
  assign _T_90405 = _T_90398[5]; // @[util.scala 33:60:@36493.4]
  assign _T_90406 = _T_90398[6]; // @[util.scala 33:60:@36494.4]
  assign _T_90407 = _T_90398[7]; // @[util.scala 33:60:@36495.4]
  assign _T_90408 = _T_90398[8]; // @[util.scala 33:60:@36496.4]
  assign _T_90409 = _T_90398[9]; // @[util.scala 33:60:@36497.4]
  assign _T_90410 = _T_90398[10]; // @[util.scala 33:60:@36498.4]
  assign _T_90411 = _T_90398[11]; // @[util.scala 33:60:@36499.4]
  assign _T_90412 = _T_90398[12]; // @[util.scala 33:60:@36500.4]
  assign _T_90413 = _T_90398[13]; // @[util.scala 33:60:@36501.4]
  assign _T_90414 = _T_90398[14]; // @[util.scala 33:60:@36502.4]
  assign _T_90415 = _T_90398[15]; // @[util.scala 33:60:@36503.4]
  assign _T_93512 = dataKnownPReg_15 == 1'h0; // @[LoadQueue.scala 229:41:@39026.4]
  assign _T_93513 = addrKnownPReg_15 & _T_93512; // @[LoadQueue.scala 229:38:@39027.4]
  assign _T_93515 = bypassInitiated_15 == 1'h0; // @[LoadQueue.scala 230:12:@39029.6]
  assign _T_93517 = prevPriorityRequest_15 == 1'h0; // @[LoadQueue.scala 230:46:@39030.6]
  assign _T_93518 = _T_93515 & _T_93517; // @[LoadQueue.scala 230:43:@39031.6]
  assign _T_93520 = dataKnown_15 == 1'h0; // @[LoadQueue.scala 230:84:@39032.6]
  assign _T_93521 = _T_93518 & _T_93520; // @[LoadQueue.scala 230:81:@39033.6]
  assign _T_93524 = storeAddrNotKnownFlagsPReg_15_0 | storeAddrNotKnownFlagsPReg_15_1; // @[LoadQueue.scala 233:86:@39036.8]
  assign _T_93525 = _T_93524 | storeAddrNotKnownFlagsPReg_15_2; // @[LoadQueue.scala 233:86:@39037.8]
  assign _T_93526 = _T_93525 | storeAddrNotKnownFlagsPReg_15_3; // @[LoadQueue.scala 233:86:@39038.8]
  assign _T_93527 = _T_93526 | storeAddrNotKnownFlagsPReg_15_4; // @[LoadQueue.scala 233:86:@39039.8]
  assign _T_93528 = _T_93527 | storeAddrNotKnownFlagsPReg_15_5; // @[LoadQueue.scala 233:86:@39040.8]
  assign _T_93529 = _T_93528 | storeAddrNotKnownFlagsPReg_15_6; // @[LoadQueue.scala 233:86:@39041.8]
  assign _T_93530 = _T_93529 | storeAddrNotKnownFlagsPReg_15_7; // @[LoadQueue.scala 233:86:@39042.8]
  assign _T_93531 = _T_93530 | storeAddrNotKnownFlagsPReg_15_8; // @[LoadQueue.scala 233:86:@39043.8]
  assign _T_93532 = _T_93531 | storeAddrNotKnownFlagsPReg_15_9; // @[LoadQueue.scala 233:86:@39044.8]
  assign _T_93533 = _T_93532 | storeAddrNotKnownFlagsPReg_15_10; // @[LoadQueue.scala 233:86:@39045.8]
  assign _T_93534 = _T_93533 | storeAddrNotKnownFlagsPReg_15_11; // @[LoadQueue.scala 233:86:@39046.8]
  assign _T_93535 = _T_93534 | storeAddrNotKnownFlagsPReg_15_12; // @[LoadQueue.scala 233:86:@39047.8]
  assign _T_93536 = _T_93535 | storeAddrNotKnownFlagsPReg_15_13; // @[LoadQueue.scala 233:86:@39048.8]
  assign _T_93537 = _T_93536 | storeAddrNotKnownFlagsPReg_15_14; // @[LoadQueue.scala 233:86:@39049.8]
  assign _T_93538 = _T_93537 | storeAddrNotKnownFlagsPReg_15_15; // @[LoadQueue.scala 233:86:@39050.8]
  assign _T_93540 = _T_93538 == 1'h0; // @[LoadQueue.scala 233:38:@39051.8]
  assign _T_93559 = _T_90338 == 1'h0; // @[LoadQueue.scala 234:11:@39068.8]
  assign _T_93560 = _T_93540 & _T_93559; // @[LoadQueue.scala 233:103:@39069.8]
  assign _GEN_2028 = _T_93521 ? _T_93560 : 1'h0; // @[LoadQueue.scala 230:110:@39034.6]
  assign loadRequest_15 = _T_93513 ? _GEN_2028 : 1'h0; // @[LoadQueue.scala 229:71:@39028.4]
  assign _T_90456 = loadRequest_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36521.4]
  assign _T_93428 = dataKnownPReg_14 == 1'h0; // @[LoadQueue.scala 229:41:@38944.4]
  assign _T_93429 = addrKnownPReg_14 & _T_93428; // @[LoadQueue.scala 229:38:@38945.4]
  assign _T_93431 = bypassInitiated_14 == 1'h0; // @[LoadQueue.scala 230:12:@38947.6]
  assign _T_93433 = prevPriorityRequest_14 == 1'h0; // @[LoadQueue.scala 230:46:@38948.6]
  assign _T_93434 = _T_93431 & _T_93433; // @[LoadQueue.scala 230:43:@38949.6]
  assign _T_93436 = dataKnown_14 == 1'h0; // @[LoadQueue.scala 230:84:@38950.6]
  assign _T_93437 = _T_93434 & _T_93436; // @[LoadQueue.scala 230:81:@38951.6]
  assign _T_93440 = storeAddrNotKnownFlagsPReg_14_0 | storeAddrNotKnownFlagsPReg_14_1; // @[LoadQueue.scala 233:86:@38954.8]
  assign _T_93441 = _T_93440 | storeAddrNotKnownFlagsPReg_14_2; // @[LoadQueue.scala 233:86:@38955.8]
  assign _T_93442 = _T_93441 | storeAddrNotKnownFlagsPReg_14_3; // @[LoadQueue.scala 233:86:@38956.8]
  assign _T_93443 = _T_93442 | storeAddrNotKnownFlagsPReg_14_4; // @[LoadQueue.scala 233:86:@38957.8]
  assign _T_93444 = _T_93443 | storeAddrNotKnownFlagsPReg_14_5; // @[LoadQueue.scala 233:86:@38958.8]
  assign _T_93445 = _T_93444 | storeAddrNotKnownFlagsPReg_14_6; // @[LoadQueue.scala 233:86:@38959.8]
  assign _T_93446 = _T_93445 | storeAddrNotKnownFlagsPReg_14_7; // @[LoadQueue.scala 233:86:@38960.8]
  assign _T_93447 = _T_93446 | storeAddrNotKnownFlagsPReg_14_8; // @[LoadQueue.scala 233:86:@38961.8]
  assign _T_93448 = _T_93447 | storeAddrNotKnownFlagsPReg_14_9; // @[LoadQueue.scala 233:86:@38962.8]
  assign _T_93449 = _T_93448 | storeAddrNotKnownFlagsPReg_14_10; // @[LoadQueue.scala 233:86:@38963.8]
  assign _T_93450 = _T_93449 | storeAddrNotKnownFlagsPReg_14_11; // @[LoadQueue.scala 233:86:@38964.8]
  assign _T_93451 = _T_93450 | storeAddrNotKnownFlagsPReg_14_12; // @[LoadQueue.scala 233:86:@38965.8]
  assign _T_93452 = _T_93451 | storeAddrNotKnownFlagsPReg_14_13; // @[LoadQueue.scala 233:86:@38966.8]
  assign _T_93453 = _T_93452 | storeAddrNotKnownFlagsPReg_14_14; // @[LoadQueue.scala 233:86:@38967.8]
  assign _T_93454 = _T_93453 | storeAddrNotKnownFlagsPReg_14_15; // @[LoadQueue.scala 233:86:@38968.8]
  assign _T_93456 = _T_93454 == 1'h0; // @[LoadQueue.scala 233:38:@38969.8]
  assign _T_93475 = _T_90202 == 1'h0; // @[LoadQueue.scala 234:11:@38986.8]
  assign _T_93476 = _T_93456 & _T_93475; // @[LoadQueue.scala 233:103:@38987.8]
  assign _GEN_2024 = _T_93437 ? _T_93476 : 1'h0; // @[LoadQueue.scala 230:110:@38952.6]
  assign loadRequest_14 = _T_93429 ? _GEN_2024 : 1'h0; // @[LoadQueue.scala 229:71:@38946.4]
  assign _T_90457 = loadRequest_14 ? 16'h4000 : _T_90456; // @[Mux.scala 31:69:@36522.4]
  assign _T_93344 = dataKnownPReg_13 == 1'h0; // @[LoadQueue.scala 229:41:@38862.4]
  assign _T_93345 = addrKnownPReg_13 & _T_93344; // @[LoadQueue.scala 229:38:@38863.4]
  assign _T_93347 = bypassInitiated_13 == 1'h0; // @[LoadQueue.scala 230:12:@38865.6]
  assign _T_93349 = prevPriorityRequest_13 == 1'h0; // @[LoadQueue.scala 230:46:@38866.6]
  assign _T_93350 = _T_93347 & _T_93349; // @[LoadQueue.scala 230:43:@38867.6]
  assign _T_93352 = dataKnown_13 == 1'h0; // @[LoadQueue.scala 230:84:@38868.6]
  assign _T_93353 = _T_93350 & _T_93352; // @[LoadQueue.scala 230:81:@38869.6]
  assign _T_93356 = storeAddrNotKnownFlagsPReg_13_0 | storeAddrNotKnownFlagsPReg_13_1; // @[LoadQueue.scala 233:86:@38872.8]
  assign _T_93357 = _T_93356 | storeAddrNotKnownFlagsPReg_13_2; // @[LoadQueue.scala 233:86:@38873.8]
  assign _T_93358 = _T_93357 | storeAddrNotKnownFlagsPReg_13_3; // @[LoadQueue.scala 233:86:@38874.8]
  assign _T_93359 = _T_93358 | storeAddrNotKnownFlagsPReg_13_4; // @[LoadQueue.scala 233:86:@38875.8]
  assign _T_93360 = _T_93359 | storeAddrNotKnownFlagsPReg_13_5; // @[LoadQueue.scala 233:86:@38876.8]
  assign _T_93361 = _T_93360 | storeAddrNotKnownFlagsPReg_13_6; // @[LoadQueue.scala 233:86:@38877.8]
  assign _T_93362 = _T_93361 | storeAddrNotKnownFlagsPReg_13_7; // @[LoadQueue.scala 233:86:@38878.8]
  assign _T_93363 = _T_93362 | storeAddrNotKnownFlagsPReg_13_8; // @[LoadQueue.scala 233:86:@38879.8]
  assign _T_93364 = _T_93363 | storeAddrNotKnownFlagsPReg_13_9; // @[LoadQueue.scala 233:86:@38880.8]
  assign _T_93365 = _T_93364 | storeAddrNotKnownFlagsPReg_13_10; // @[LoadQueue.scala 233:86:@38881.8]
  assign _T_93366 = _T_93365 | storeAddrNotKnownFlagsPReg_13_11; // @[LoadQueue.scala 233:86:@38882.8]
  assign _T_93367 = _T_93366 | storeAddrNotKnownFlagsPReg_13_12; // @[LoadQueue.scala 233:86:@38883.8]
  assign _T_93368 = _T_93367 | storeAddrNotKnownFlagsPReg_13_13; // @[LoadQueue.scala 233:86:@38884.8]
  assign _T_93369 = _T_93368 | storeAddrNotKnownFlagsPReg_13_14; // @[LoadQueue.scala 233:86:@38885.8]
  assign _T_93370 = _T_93369 | storeAddrNotKnownFlagsPReg_13_15; // @[LoadQueue.scala 233:86:@38886.8]
  assign _T_93372 = _T_93370 == 1'h0; // @[LoadQueue.scala 233:38:@38887.8]
  assign _T_93391 = _T_90066 == 1'h0; // @[LoadQueue.scala 234:11:@38904.8]
  assign _T_93392 = _T_93372 & _T_93391; // @[LoadQueue.scala 233:103:@38905.8]
  assign _GEN_2020 = _T_93353 ? _T_93392 : 1'h0; // @[LoadQueue.scala 230:110:@38870.6]
  assign loadRequest_13 = _T_93345 ? _GEN_2020 : 1'h0; // @[LoadQueue.scala 229:71:@38864.4]
  assign _T_90458 = loadRequest_13 ? 16'h2000 : _T_90457; // @[Mux.scala 31:69:@36523.4]
  assign _T_93260 = dataKnownPReg_12 == 1'h0; // @[LoadQueue.scala 229:41:@38780.4]
  assign _T_93261 = addrKnownPReg_12 & _T_93260; // @[LoadQueue.scala 229:38:@38781.4]
  assign _T_93263 = bypassInitiated_12 == 1'h0; // @[LoadQueue.scala 230:12:@38783.6]
  assign _T_93265 = prevPriorityRequest_12 == 1'h0; // @[LoadQueue.scala 230:46:@38784.6]
  assign _T_93266 = _T_93263 & _T_93265; // @[LoadQueue.scala 230:43:@38785.6]
  assign _T_93268 = dataKnown_12 == 1'h0; // @[LoadQueue.scala 230:84:@38786.6]
  assign _T_93269 = _T_93266 & _T_93268; // @[LoadQueue.scala 230:81:@38787.6]
  assign _T_93272 = storeAddrNotKnownFlagsPReg_12_0 | storeAddrNotKnownFlagsPReg_12_1; // @[LoadQueue.scala 233:86:@38790.8]
  assign _T_93273 = _T_93272 | storeAddrNotKnownFlagsPReg_12_2; // @[LoadQueue.scala 233:86:@38791.8]
  assign _T_93274 = _T_93273 | storeAddrNotKnownFlagsPReg_12_3; // @[LoadQueue.scala 233:86:@38792.8]
  assign _T_93275 = _T_93274 | storeAddrNotKnownFlagsPReg_12_4; // @[LoadQueue.scala 233:86:@38793.8]
  assign _T_93276 = _T_93275 | storeAddrNotKnownFlagsPReg_12_5; // @[LoadQueue.scala 233:86:@38794.8]
  assign _T_93277 = _T_93276 | storeAddrNotKnownFlagsPReg_12_6; // @[LoadQueue.scala 233:86:@38795.8]
  assign _T_93278 = _T_93277 | storeAddrNotKnownFlagsPReg_12_7; // @[LoadQueue.scala 233:86:@38796.8]
  assign _T_93279 = _T_93278 | storeAddrNotKnownFlagsPReg_12_8; // @[LoadQueue.scala 233:86:@38797.8]
  assign _T_93280 = _T_93279 | storeAddrNotKnownFlagsPReg_12_9; // @[LoadQueue.scala 233:86:@38798.8]
  assign _T_93281 = _T_93280 | storeAddrNotKnownFlagsPReg_12_10; // @[LoadQueue.scala 233:86:@38799.8]
  assign _T_93282 = _T_93281 | storeAddrNotKnownFlagsPReg_12_11; // @[LoadQueue.scala 233:86:@38800.8]
  assign _T_93283 = _T_93282 | storeAddrNotKnownFlagsPReg_12_12; // @[LoadQueue.scala 233:86:@38801.8]
  assign _T_93284 = _T_93283 | storeAddrNotKnownFlagsPReg_12_13; // @[LoadQueue.scala 233:86:@38802.8]
  assign _T_93285 = _T_93284 | storeAddrNotKnownFlagsPReg_12_14; // @[LoadQueue.scala 233:86:@38803.8]
  assign _T_93286 = _T_93285 | storeAddrNotKnownFlagsPReg_12_15; // @[LoadQueue.scala 233:86:@38804.8]
  assign _T_93288 = _T_93286 == 1'h0; // @[LoadQueue.scala 233:38:@38805.8]
  assign _T_93307 = _T_89930 == 1'h0; // @[LoadQueue.scala 234:11:@38822.8]
  assign _T_93308 = _T_93288 & _T_93307; // @[LoadQueue.scala 233:103:@38823.8]
  assign _GEN_2016 = _T_93269 ? _T_93308 : 1'h0; // @[LoadQueue.scala 230:110:@38788.6]
  assign loadRequest_12 = _T_93261 ? _GEN_2016 : 1'h0; // @[LoadQueue.scala 229:71:@38782.4]
  assign _T_90459 = loadRequest_12 ? 16'h1000 : _T_90458; // @[Mux.scala 31:69:@36524.4]
  assign _T_93176 = dataKnownPReg_11 == 1'h0; // @[LoadQueue.scala 229:41:@38698.4]
  assign _T_93177 = addrKnownPReg_11 & _T_93176; // @[LoadQueue.scala 229:38:@38699.4]
  assign _T_93179 = bypassInitiated_11 == 1'h0; // @[LoadQueue.scala 230:12:@38701.6]
  assign _T_93181 = prevPriorityRequest_11 == 1'h0; // @[LoadQueue.scala 230:46:@38702.6]
  assign _T_93182 = _T_93179 & _T_93181; // @[LoadQueue.scala 230:43:@38703.6]
  assign _T_93184 = dataKnown_11 == 1'h0; // @[LoadQueue.scala 230:84:@38704.6]
  assign _T_93185 = _T_93182 & _T_93184; // @[LoadQueue.scala 230:81:@38705.6]
  assign _T_93188 = storeAddrNotKnownFlagsPReg_11_0 | storeAddrNotKnownFlagsPReg_11_1; // @[LoadQueue.scala 233:86:@38708.8]
  assign _T_93189 = _T_93188 | storeAddrNotKnownFlagsPReg_11_2; // @[LoadQueue.scala 233:86:@38709.8]
  assign _T_93190 = _T_93189 | storeAddrNotKnownFlagsPReg_11_3; // @[LoadQueue.scala 233:86:@38710.8]
  assign _T_93191 = _T_93190 | storeAddrNotKnownFlagsPReg_11_4; // @[LoadQueue.scala 233:86:@38711.8]
  assign _T_93192 = _T_93191 | storeAddrNotKnownFlagsPReg_11_5; // @[LoadQueue.scala 233:86:@38712.8]
  assign _T_93193 = _T_93192 | storeAddrNotKnownFlagsPReg_11_6; // @[LoadQueue.scala 233:86:@38713.8]
  assign _T_93194 = _T_93193 | storeAddrNotKnownFlagsPReg_11_7; // @[LoadQueue.scala 233:86:@38714.8]
  assign _T_93195 = _T_93194 | storeAddrNotKnownFlagsPReg_11_8; // @[LoadQueue.scala 233:86:@38715.8]
  assign _T_93196 = _T_93195 | storeAddrNotKnownFlagsPReg_11_9; // @[LoadQueue.scala 233:86:@38716.8]
  assign _T_93197 = _T_93196 | storeAddrNotKnownFlagsPReg_11_10; // @[LoadQueue.scala 233:86:@38717.8]
  assign _T_93198 = _T_93197 | storeAddrNotKnownFlagsPReg_11_11; // @[LoadQueue.scala 233:86:@38718.8]
  assign _T_93199 = _T_93198 | storeAddrNotKnownFlagsPReg_11_12; // @[LoadQueue.scala 233:86:@38719.8]
  assign _T_93200 = _T_93199 | storeAddrNotKnownFlagsPReg_11_13; // @[LoadQueue.scala 233:86:@38720.8]
  assign _T_93201 = _T_93200 | storeAddrNotKnownFlagsPReg_11_14; // @[LoadQueue.scala 233:86:@38721.8]
  assign _T_93202 = _T_93201 | storeAddrNotKnownFlagsPReg_11_15; // @[LoadQueue.scala 233:86:@38722.8]
  assign _T_93204 = _T_93202 == 1'h0; // @[LoadQueue.scala 233:38:@38723.8]
  assign _T_93223 = _T_89794 == 1'h0; // @[LoadQueue.scala 234:11:@38740.8]
  assign _T_93224 = _T_93204 & _T_93223; // @[LoadQueue.scala 233:103:@38741.8]
  assign _GEN_2012 = _T_93185 ? _T_93224 : 1'h0; // @[LoadQueue.scala 230:110:@38706.6]
  assign loadRequest_11 = _T_93177 ? _GEN_2012 : 1'h0; // @[LoadQueue.scala 229:71:@38700.4]
  assign _T_90460 = loadRequest_11 ? 16'h800 : _T_90459; // @[Mux.scala 31:69:@36525.4]
  assign _T_93092 = dataKnownPReg_10 == 1'h0; // @[LoadQueue.scala 229:41:@38616.4]
  assign _T_93093 = addrKnownPReg_10 & _T_93092; // @[LoadQueue.scala 229:38:@38617.4]
  assign _T_93095 = bypassInitiated_10 == 1'h0; // @[LoadQueue.scala 230:12:@38619.6]
  assign _T_93097 = prevPriorityRequest_10 == 1'h0; // @[LoadQueue.scala 230:46:@38620.6]
  assign _T_93098 = _T_93095 & _T_93097; // @[LoadQueue.scala 230:43:@38621.6]
  assign _T_93100 = dataKnown_10 == 1'h0; // @[LoadQueue.scala 230:84:@38622.6]
  assign _T_93101 = _T_93098 & _T_93100; // @[LoadQueue.scala 230:81:@38623.6]
  assign _T_93104 = storeAddrNotKnownFlagsPReg_10_0 | storeAddrNotKnownFlagsPReg_10_1; // @[LoadQueue.scala 233:86:@38626.8]
  assign _T_93105 = _T_93104 | storeAddrNotKnownFlagsPReg_10_2; // @[LoadQueue.scala 233:86:@38627.8]
  assign _T_93106 = _T_93105 | storeAddrNotKnownFlagsPReg_10_3; // @[LoadQueue.scala 233:86:@38628.8]
  assign _T_93107 = _T_93106 | storeAddrNotKnownFlagsPReg_10_4; // @[LoadQueue.scala 233:86:@38629.8]
  assign _T_93108 = _T_93107 | storeAddrNotKnownFlagsPReg_10_5; // @[LoadQueue.scala 233:86:@38630.8]
  assign _T_93109 = _T_93108 | storeAddrNotKnownFlagsPReg_10_6; // @[LoadQueue.scala 233:86:@38631.8]
  assign _T_93110 = _T_93109 | storeAddrNotKnownFlagsPReg_10_7; // @[LoadQueue.scala 233:86:@38632.8]
  assign _T_93111 = _T_93110 | storeAddrNotKnownFlagsPReg_10_8; // @[LoadQueue.scala 233:86:@38633.8]
  assign _T_93112 = _T_93111 | storeAddrNotKnownFlagsPReg_10_9; // @[LoadQueue.scala 233:86:@38634.8]
  assign _T_93113 = _T_93112 | storeAddrNotKnownFlagsPReg_10_10; // @[LoadQueue.scala 233:86:@38635.8]
  assign _T_93114 = _T_93113 | storeAddrNotKnownFlagsPReg_10_11; // @[LoadQueue.scala 233:86:@38636.8]
  assign _T_93115 = _T_93114 | storeAddrNotKnownFlagsPReg_10_12; // @[LoadQueue.scala 233:86:@38637.8]
  assign _T_93116 = _T_93115 | storeAddrNotKnownFlagsPReg_10_13; // @[LoadQueue.scala 233:86:@38638.8]
  assign _T_93117 = _T_93116 | storeAddrNotKnownFlagsPReg_10_14; // @[LoadQueue.scala 233:86:@38639.8]
  assign _T_93118 = _T_93117 | storeAddrNotKnownFlagsPReg_10_15; // @[LoadQueue.scala 233:86:@38640.8]
  assign _T_93120 = _T_93118 == 1'h0; // @[LoadQueue.scala 233:38:@38641.8]
  assign _T_93139 = _T_89658 == 1'h0; // @[LoadQueue.scala 234:11:@38658.8]
  assign _T_93140 = _T_93120 & _T_93139; // @[LoadQueue.scala 233:103:@38659.8]
  assign _GEN_2008 = _T_93101 ? _T_93140 : 1'h0; // @[LoadQueue.scala 230:110:@38624.6]
  assign loadRequest_10 = _T_93093 ? _GEN_2008 : 1'h0; // @[LoadQueue.scala 229:71:@38618.4]
  assign _T_90461 = loadRequest_10 ? 16'h400 : _T_90460; // @[Mux.scala 31:69:@36526.4]
  assign _T_93008 = dataKnownPReg_9 == 1'h0; // @[LoadQueue.scala 229:41:@38534.4]
  assign _T_93009 = addrKnownPReg_9 & _T_93008; // @[LoadQueue.scala 229:38:@38535.4]
  assign _T_93011 = bypassInitiated_9 == 1'h0; // @[LoadQueue.scala 230:12:@38537.6]
  assign _T_93013 = prevPriorityRequest_9 == 1'h0; // @[LoadQueue.scala 230:46:@38538.6]
  assign _T_93014 = _T_93011 & _T_93013; // @[LoadQueue.scala 230:43:@38539.6]
  assign _T_93016 = dataKnown_9 == 1'h0; // @[LoadQueue.scala 230:84:@38540.6]
  assign _T_93017 = _T_93014 & _T_93016; // @[LoadQueue.scala 230:81:@38541.6]
  assign _T_93020 = storeAddrNotKnownFlagsPReg_9_0 | storeAddrNotKnownFlagsPReg_9_1; // @[LoadQueue.scala 233:86:@38544.8]
  assign _T_93021 = _T_93020 | storeAddrNotKnownFlagsPReg_9_2; // @[LoadQueue.scala 233:86:@38545.8]
  assign _T_93022 = _T_93021 | storeAddrNotKnownFlagsPReg_9_3; // @[LoadQueue.scala 233:86:@38546.8]
  assign _T_93023 = _T_93022 | storeAddrNotKnownFlagsPReg_9_4; // @[LoadQueue.scala 233:86:@38547.8]
  assign _T_93024 = _T_93023 | storeAddrNotKnownFlagsPReg_9_5; // @[LoadQueue.scala 233:86:@38548.8]
  assign _T_93025 = _T_93024 | storeAddrNotKnownFlagsPReg_9_6; // @[LoadQueue.scala 233:86:@38549.8]
  assign _T_93026 = _T_93025 | storeAddrNotKnownFlagsPReg_9_7; // @[LoadQueue.scala 233:86:@38550.8]
  assign _T_93027 = _T_93026 | storeAddrNotKnownFlagsPReg_9_8; // @[LoadQueue.scala 233:86:@38551.8]
  assign _T_93028 = _T_93027 | storeAddrNotKnownFlagsPReg_9_9; // @[LoadQueue.scala 233:86:@38552.8]
  assign _T_93029 = _T_93028 | storeAddrNotKnownFlagsPReg_9_10; // @[LoadQueue.scala 233:86:@38553.8]
  assign _T_93030 = _T_93029 | storeAddrNotKnownFlagsPReg_9_11; // @[LoadQueue.scala 233:86:@38554.8]
  assign _T_93031 = _T_93030 | storeAddrNotKnownFlagsPReg_9_12; // @[LoadQueue.scala 233:86:@38555.8]
  assign _T_93032 = _T_93031 | storeAddrNotKnownFlagsPReg_9_13; // @[LoadQueue.scala 233:86:@38556.8]
  assign _T_93033 = _T_93032 | storeAddrNotKnownFlagsPReg_9_14; // @[LoadQueue.scala 233:86:@38557.8]
  assign _T_93034 = _T_93033 | storeAddrNotKnownFlagsPReg_9_15; // @[LoadQueue.scala 233:86:@38558.8]
  assign _T_93036 = _T_93034 == 1'h0; // @[LoadQueue.scala 233:38:@38559.8]
  assign _T_93055 = _T_89522 == 1'h0; // @[LoadQueue.scala 234:11:@38576.8]
  assign _T_93056 = _T_93036 & _T_93055; // @[LoadQueue.scala 233:103:@38577.8]
  assign _GEN_2004 = _T_93017 ? _T_93056 : 1'h0; // @[LoadQueue.scala 230:110:@38542.6]
  assign loadRequest_9 = _T_93009 ? _GEN_2004 : 1'h0; // @[LoadQueue.scala 229:71:@38536.4]
  assign _T_90462 = loadRequest_9 ? 16'h200 : _T_90461; // @[Mux.scala 31:69:@36527.4]
  assign _T_92924 = dataKnownPReg_8 == 1'h0; // @[LoadQueue.scala 229:41:@38452.4]
  assign _T_92925 = addrKnownPReg_8 & _T_92924; // @[LoadQueue.scala 229:38:@38453.4]
  assign _T_92927 = bypassInitiated_8 == 1'h0; // @[LoadQueue.scala 230:12:@38455.6]
  assign _T_92929 = prevPriorityRequest_8 == 1'h0; // @[LoadQueue.scala 230:46:@38456.6]
  assign _T_92930 = _T_92927 & _T_92929; // @[LoadQueue.scala 230:43:@38457.6]
  assign _T_92932 = dataKnown_8 == 1'h0; // @[LoadQueue.scala 230:84:@38458.6]
  assign _T_92933 = _T_92930 & _T_92932; // @[LoadQueue.scala 230:81:@38459.6]
  assign _T_92936 = storeAddrNotKnownFlagsPReg_8_0 | storeAddrNotKnownFlagsPReg_8_1; // @[LoadQueue.scala 233:86:@38462.8]
  assign _T_92937 = _T_92936 | storeAddrNotKnownFlagsPReg_8_2; // @[LoadQueue.scala 233:86:@38463.8]
  assign _T_92938 = _T_92937 | storeAddrNotKnownFlagsPReg_8_3; // @[LoadQueue.scala 233:86:@38464.8]
  assign _T_92939 = _T_92938 | storeAddrNotKnownFlagsPReg_8_4; // @[LoadQueue.scala 233:86:@38465.8]
  assign _T_92940 = _T_92939 | storeAddrNotKnownFlagsPReg_8_5; // @[LoadQueue.scala 233:86:@38466.8]
  assign _T_92941 = _T_92940 | storeAddrNotKnownFlagsPReg_8_6; // @[LoadQueue.scala 233:86:@38467.8]
  assign _T_92942 = _T_92941 | storeAddrNotKnownFlagsPReg_8_7; // @[LoadQueue.scala 233:86:@38468.8]
  assign _T_92943 = _T_92942 | storeAddrNotKnownFlagsPReg_8_8; // @[LoadQueue.scala 233:86:@38469.8]
  assign _T_92944 = _T_92943 | storeAddrNotKnownFlagsPReg_8_9; // @[LoadQueue.scala 233:86:@38470.8]
  assign _T_92945 = _T_92944 | storeAddrNotKnownFlagsPReg_8_10; // @[LoadQueue.scala 233:86:@38471.8]
  assign _T_92946 = _T_92945 | storeAddrNotKnownFlagsPReg_8_11; // @[LoadQueue.scala 233:86:@38472.8]
  assign _T_92947 = _T_92946 | storeAddrNotKnownFlagsPReg_8_12; // @[LoadQueue.scala 233:86:@38473.8]
  assign _T_92948 = _T_92947 | storeAddrNotKnownFlagsPReg_8_13; // @[LoadQueue.scala 233:86:@38474.8]
  assign _T_92949 = _T_92948 | storeAddrNotKnownFlagsPReg_8_14; // @[LoadQueue.scala 233:86:@38475.8]
  assign _T_92950 = _T_92949 | storeAddrNotKnownFlagsPReg_8_15; // @[LoadQueue.scala 233:86:@38476.8]
  assign _T_92952 = _T_92950 == 1'h0; // @[LoadQueue.scala 233:38:@38477.8]
  assign _T_92971 = _T_89386 == 1'h0; // @[LoadQueue.scala 234:11:@38494.8]
  assign _T_92972 = _T_92952 & _T_92971; // @[LoadQueue.scala 233:103:@38495.8]
  assign _GEN_2000 = _T_92933 ? _T_92972 : 1'h0; // @[LoadQueue.scala 230:110:@38460.6]
  assign loadRequest_8 = _T_92925 ? _GEN_2000 : 1'h0; // @[LoadQueue.scala 229:71:@38454.4]
  assign _T_90463 = loadRequest_8 ? 16'h100 : _T_90462; // @[Mux.scala 31:69:@36528.4]
  assign _T_92840 = dataKnownPReg_7 == 1'h0; // @[LoadQueue.scala 229:41:@38370.4]
  assign _T_92841 = addrKnownPReg_7 & _T_92840; // @[LoadQueue.scala 229:38:@38371.4]
  assign _T_92843 = bypassInitiated_7 == 1'h0; // @[LoadQueue.scala 230:12:@38373.6]
  assign _T_92845 = prevPriorityRequest_7 == 1'h0; // @[LoadQueue.scala 230:46:@38374.6]
  assign _T_92846 = _T_92843 & _T_92845; // @[LoadQueue.scala 230:43:@38375.6]
  assign _T_92848 = dataKnown_7 == 1'h0; // @[LoadQueue.scala 230:84:@38376.6]
  assign _T_92849 = _T_92846 & _T_92848; // @[LoadQueue.scala 230:81:@38377.6]
  assign _T_92852 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[LoadQueue.scala 233:86:@38380.8]
  assign _T_92853 = _T_92852 | storeAddrNotKnownFlagsPReg_7_2; // @[LoadQueue.scala 233:86:@38381.8]
  assign _T_92854 = _T_92853 | storeAddrNotKnownFlagsPReg_7_3; // @[LoadQueue.scala 233:86:@38382.8]
  assign _T_92855 = _T_92854 | storeAddrNotKnownFlagsPReg_7_4; // @[LoadQueue.scala 233:86:@38383.8]
  assign _T_92856 = _T_92855 | storeAddrNotKnownFlagsPReg_7_5; // @[LoadQueue.scala 233:86:@38384.8]
  assign _T_92857 = _T_92856 | storeAddrNotKnownFlagsPReg_7_6; // @[LoadQueue.scala 233:86:@38385.8]
  assign _T_92858 = _T_92857 | storeAddrNotKnownFlagsPReg_7_7; // @[LoadQueue.scala 233:86:@38386.8]
  assign _T_92859 = _T_92858 | storeAddrNotKnownFlagsPReg_7_8; // @[LoadQueue.scala 233:86:@38387.8]
  assign _T_92860 = _T_92859 | storeAddrNotKnownFlagsPReg_7_9; // @[LoadQueue.scala 233:86:@38388.8]
  assign _T_92861 = _T_92860 | storeAddrNotKnownFlagsPReg_7_10; // @[LoadQueue.scala 233:86:@38389.8]
  assign _T_92862 = _T_92861 | storeAddrNotKnownFlagsPReg_7_11; // @[LoadQueue.scala 233:86:@38390.8]
  assign _T_92863 = _T_92862 | storeAddrNotKnownFlagsPReg_7_12; // @[LoadQueue.scala 233:86:@38391.8]
  assign _T_92864 = _T_92863 | storeAddrNotKnownFlagsPReg_7_13; // @[LoadQueue.scala 233:86:@38392.8]
  assign _T_92865 = _T_92864 | storeAddrNotKnownFlagsPReg_7_14; // @[LoadQueue.scala 233:86:@38393.8]
  assign _T_92866 = _T_92865 | storeAddrNotKnownFlagsPReg_7_15; // @[LoadQueue.scala 233:86:@38394.8]
  assign _T_92868 = _T_92866 == 1'h0; // @[LoadQueue.scala 233:38:@38395.8]
  assign _T_92887 = _T_89250 == 1'h0; // @[LoadQueue.scala 234:11:@38412.8]
  assign _T_92888 = _T_92868 & _T_92887; // @[LoadQueue.scala 233:103:@38413.8]
  assign _GEN_1996 = _T_92849 ? _T_92888 : 1'h0; // @[LoadQueue.scala 230:110:@38378.6]
  assign loadRequest_7 = _T_92841 ? _GEN_1996 : 1'h0; // @[LoadQueue.scala 229:71:@38372.4]
  assign _T_90464 = loadRequest_7 ? 16'h80 : _T_90463; // @[Mux.scala 31:69:@36529.4]
  assign _T_92756 = dataKnownPReg_6 == 1'h0; // @[LoadQueue.scala 229:41:@38288.4]
  assign _T_92757 = addrKnownPReg_6 & _T_92756; // @[LoadQueue.scala 229:38:@38289.4]
  assign _T_92759 = bypassInitiated_6 == 1'h0; // @[LoadQueue.scala 230:12:@38291.6]
  assign _T_92761 = prevPriorityRequest_6 == 1'h0; // @[LoadQueue.scala 230:46:@38292.6]
  assign _T_92762 = _T_92759 & _T_92761; // @[LoadQueue.scala 230:43:@38293.6]
  assign _T_92764 = dataKnown_6 == 1'h0; // @[LoadQueue.scala 230:84:@38294.6]
  assign _T_92765 = _T_92762 & _T_92764; // @[LoadQueue.scala 230:81:@38295.6]
  assign _T_92768 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[LoadQueue.scala 233:86:@38298.8]
  assign _T_92769 = _T_92768 | storeAddrNotKnownFlagsPReg_6_2; // @[LoadQueue.scala 233:86:@38299.8]
  assign _T_92770 = _T_92769 | storeAddrNotKnownFlagsPReg_6_3; // @[LoadQueue.scala 233:86:@38300.8]
  assign _T_92771 = _T_92770 | storeAddrNotKnownFlagsPReg_6_4; // @[LoadQueue.scala 233:86:@38301.8]
  assign _T_92772 = _T_92771 | storeAddrNotKnownFlagsPReg_6_5; // @[LoadQueue.scala 233:86:@38302.8]
  assign _T_92773 = _T_92772 | storeAddrNotKnownFlagsPReg_6_6; // @[LoadQueue.scala 233:86:@38303.8]
  assign _T_92774 = _T_92773 | storeAddrNotKnownFlagsPReg_6_7; // @[LoadQueue.scala 233:86:@38304.8]
  assign _T_92775 = _T_92774 | storeAddrNotKnownFlagsPReg_6_8; // @[LoadQueue.scala 233:86:@38305.8]
  assign _T_92776 = _T_92775 | storeAddrNotKnownFlagsPReg_6_9; // @[LoadQueue.scala 233:86:@38306.8]
  assign _T_92777 = _T_92776 | storeAddrNotKnownFlagsPReg_6_10; // @[LoadQueue.scala 233:86:@38307.8]
  assign _T_92778 = _T_92777 | storeAddrNotKnownFlagsPReg_6_11; // @[LoadQueue.scala 233:86:@38308.8]
  assign _T_92779 = _T_92778 | storeAddrNotKnownFlagsPReg_6_12; // @[LoadQueue.scala 233:86:@38309.8]
  assign _T_92780 = _T_92779 | storeAddrNotKnownFlagsPReg_6_13; // @[LoadQueue.scala 233:86:@38310.8]
  assign _T_92781 = _T_92780 | storeAddrNotKnownFlagsPReg_6_14; // @[LoadQueue.scala 233:86:@38311.8]
  assign _T_92782 = _T_92781 | storeAddrNotKnownFlagsPReg_6_15; // @[LoadQueue.scala 233:86:@38312.8]
  assign _T_92784 = _T_92782 == 1'h0; // @[LoadQueue.scala 233:38:@38313.8]
  assign _T_92803 = _T_89114 == 1'h0; // @[LoadQueue.scala 234:11:@38330.8]
  assign _T_92804 = _T_92784 & _T_92803; // @[LoadQueue.scala 233:103:@38331.8]
  assign _GEN_1992 = _T_92765 ? _T_92804 : 1'h0; // @[LoadQueue.scala 230:110:@38296.6]
  assign loadRequest_6 = _T_92757 ? _GEN_1992 : 1'h0; // @[LoadQueue.scala 229:71:@38290.4]
  assign _T_90465 = loadRequest_6 ? 16'h40 : _T_90464; // @[Mux.scala 31:69:@36530.4]
  assign _T_92672 = dataKnownPReg_5 == 1'h0; // @[LoadQueue.scala 229:41:@38206.4]
  assign _T_92673 = addrKnownPReg_5 & _T_92672; // @[LoadQueue.scala 229:38:@38207.4]
  assign _T_92675 = bypassInitiated_5 == 1'h0; // @[LoadQueue.scala 230:12:@38209.6]
  assign _T_92677 = prevPriorityRequest_5 == 1'h0; // @[LoadQueue.scala 230:46:@38210.6]
  assign _T_92678 = _T_92675 & _T_92677; // @[LoadQueue.scala 230:43:@38211.6]
  assign _T_92680 = dataKnown_5 == 1'h0; // @[LoadQueue.scala 230:84:@38212.6]
  assign _T_92681 = _T_92678 & _T_92680; // @[LoadQueue.scala 230:81:@38213.6]
  assign _T_92684 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[LoadQueue.scala 233:86:@38216.8]
  assign _T_92685 = _T_92684 | storeAddrNotKnownFlagsPReg_5_2; // @[LoadQueue.scala 233:86:@38217.8]
  assign _T_92686 = _T_92685 | storeAddrNotKnownFlagsPReg_5_3; // @[LoadQueue.scala 233:86:@38218.8]
  assign _T_92687 = _T_92686 | storeAddrNotKnownFlagsPReg_5_4; // @[LoadQueue.scala 233:86:@38219.8]
  assign _T_92688 = _T_92687 | storeAddrNotKnownFlagsPReg_5_5; // @[LoadQueue.scala 233:86:@38220.8]
  assign _T_92689 = _T_92688 | storeAddrNotKnownFlagsPReg_5_6; // @[LoadQueue.scala 233:86:@38221.8]
  assign _T_92690 = _T_92689 | storeAddrNotKnownFlagsPReg_5_7; // @[LoadQueue.scala 233:86:@38222.8]
  assign _T_92691 = _T_92690 | storeAddrNotKnownFlagsPReg_5_8; // @[LoadQueue.scala 233:86:@38223.8]
  assign _T_92692 = _T_92691 | storeAddrNotKnownFlagsPReg_5_9; // @[LoadQueue.scala 233:86:@38224.8]
  assign _T_92693 = _T_92692 | storeAddrNotKnownFlagsPReg_5_10; // @[LoadQueue.scala 233:86:@38225.8]
  assign _T_92694 = _T_92693 | storeAddrNotKnownFlagsPReg_5_11; // @[LoadQueue.scala 233:86:@38226.8]
  assign _T_92695 = _T_92694 | storeAddrNotKnownFlagsPReg_5_12; // @[LoadQueue.scala 233:86:@38227.8]
  assign _T_92696 = _T_92695 | storeAddrNotKnownFlagsPReg_5_13; // @[LoadQueue.scala 233:86:@38228.8]
  assign _T_92697 = _T_92696 | storeAddrNotKnownFlagsPReg_5_14; // @[LoadQueue.scala 233:86:@38229.8]
  assign _T_92698 = _T_92697 | storeAddrNotKnownFlagsPReg_5_15; // @[LoadQueue.scala 233:86:@38230.8]
  assign _T_92700 = _T_92698 == 1'h0; // @[LoadQueue.scala 233:38:@38231.8]
  assign _T_92719 = _T_88978 == 1'h0; // @[LoadQueue.scala 234:11:@38248.8]
  assign _T_92720 = _T_92700 & _T_92719; // @[LoadQueue.scala 233:103:@38249.8]
  assign _GEN_1988 = _T_92681 ? _T_92720 : 1'h0; // @[LoadQueue.scala 230:110:@38214.6]
  assign loadRequest_5 = _T_92673 ? _GEN_1988 : 1'h0; // @[LoadQueue.scala 229:71:@38208.4]
  assign _T_90466 = loadRequest_5 ? 16'h20 : _T_90465; // @[Mux.scala 31:69:@36531.4]
  assign _T_92588 = dataKnownPReg_4 == 1'h0; // @[LoadQueue.scala 229:41:@38124.4]
  assign _T_92589 = addrKnownPReg_4 & _T_92588; // @[LoadQueue.scala 229:38:@38125.4]
  assign _T_92591 = bypassInitiated_4 == 1'h0; // @[LoadQueue.scala 230:12:@38127.6]
  assign _T_92593 = prevPriorityRequest_4 == 1'h0; // @[LoadQueue.scala 230:46:@38128.6]
  assign _T_92594 = _T_92591 & _T_92593; // @[LoadQueue.scala 230:43:@38129.6]
  assign _T_92596 = dataKnown_4 == 1'h0; // @[LoadQueue.scala 230:84:@38130.6]
  assign _T_92597 = _T_92594 & _T_92596; // @[LoadQueue.scala 230:81:@38131.6]
  assign _T_92600 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[LoadQueue.scala 233:86:@38134.8]
  assign _T_92601 = _T_92600 | storeAddrNotKnownFlagsPReg_4_2; // @[LoadQueue.scala 233:86:@38135.8]
  assign _T_92602 = _T_92601 | storeAddrNotKnownFlagsPReg_4_3; // @[LoadQueue.scala 233:86:@38136.8]
  assign _T_92603 = _T_92602 | storeAddrNotKnownFlagsPReg_4_4; // @[LoadQueue.scala 233:86:@38137.8]
  assign _T_92604 = _T_92603 | storeAddrNotKnownFlagsPReg_4_5; // @[LoadQueue.scala 233:86:@38138.8]
  assign _T_92605 = _T_92604 | storeAddrNotKnownFlagsPReg_4_6; // @[LoadQueue.scala 233:86:@38139.8]
  assign _T_92606 = _T_92605 | storeAddrNotKnownFlagsPReg_4_7; // @[LoadQueue.scala 233:86:@38140.8]
  assign _T_92607 = _T_92606 | storeAddrNotKnownFlagsPReg_4_8; // @[LoadQueue.scala 233:86:@38141.8]
  assign _T_92608 = _T_92607 | storeAddrNotKnownFlagsPReg_4_9; // @[LoadQueue.scala 233:86:@38142.8]
  assign _T_92609 = _T_92608 | storeAddrNotKnownFlagsPReg_4_10; // @[LoadQueue.scala 233:86:@38143.8]
  assign _T_92610 = _T_92609 | storeAddrNotKnownFlagsPReg_4_11; // @[LoadQueue.scala 233:86:@38144.8]
  assign _T_92611 = _T_92610 | storeAddrNotKnownFlagsPReg_4_12; // @[LoadQueue.scala 233:86:@38145.8]
  assign _T_92612 = _T_92611 | storeAddrNotKnownFlagsPReg_4_13; // @[LoadQueue.scala 233:86:@38146.8]
  assign _T_92613 = _T_92612 | storeAddrNotKnownFlagsPReg_4_14; // @[LoadQueue.scala 233:86:@38147.8]
  assign _T_92614 = _T_92613 | storeAddrNotKnownFlagsPReg_4_15; // @[LoadQueue.scala 233:86:@38148.8]
  assign _T_92616 = _T_92614 == 1'h0; // @[LoadQueue.scala 233:38:@38149.8]
  assign _T_92635 = _T_88842 == 1'h0; // @[LoadQueue.scala 234:11:@38166.8]
  assign _T_92636 = _T_92616 & _T_92635; // @[LoadQueue.scala 233:103:@38167.8]
  assign _GEN_1984 = _T_92597 ? _T_92636 : 1'h0; // @[LoadQueue.scala 230:110:@38132.6]
  assign loadRequest_4 = _T_92589 ? _GEN_1984 : 1'h0; // @[LoadQueue.scala 229:71:@38126.4]
  assign _T_90467 = loadRequest_4 ? 16'h10 : _T_90466; // @[Mux.scala 31:69:@36532.4]
  assign _T_92504 = dataKnownPReg_3 == 1'h0; // @[LoadQueue.scala 229:41:@38042.4]
  assign _T_92505 = addrKnownPReg_3 & _T_92504; // @[LoadQueue.scala 229:38:@38043.4]
  assign _T_92507 = bypassInitiated_3 == 1'h0; // @[LoadQueue.scala 230:12:@38045.6]
  assign _T_92509 = prevPriorityRequest_3 == 1'h0; // @[LoadQueue.scala 230:46:@38046.6]
  assign _T_92510 = _T_92507 & _T_92509; // @[LoadQueue.scala 230:43:@38047.6]
  assign _T_92512 = dataKnown_3 == 1'h0; // @[LoadQueue.scala 230:84:@38048.6]
  assign _T_92513 = _T_92510 & _T_92512; // @[LoadQueue.scala 230:81:@38049.6]
  assign _T_92516 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[LoadQueue.scala 233:86:@38052.8]
  assign _T_92517 = _T_92516 | storeAddrNotKnownFlagsPReg_3_2; // @[LoadQueue.scala 233:86:@38053.8]
  assign _T_92518 = _T_92517 | storeAddrNotKnownFlagsPReg_3_3; // @[LoadQueue.scala 233:86:@38054.8]
  assign _T_92519 = _T_92518 | storeAddrNotKnownFlagsPReg_3_4; // @[LoadQueue.scala 233:86:@38055.8]
  assign _T_92520 = _T_92519 | storeAddrNotKnownFlagsPReg_3_5; // @[LoadQueue.scala 233:86:@38056.8]
  assign _T_92521 = _T_92520 | storeAddrNotKnownFlagsPReg_3_6; // @[LoadQueue.scala 233:86:@38057.8]
  assign _T_92522 = _T_92521 | storeAddrNotKnownFlagsPReg_3_7; // @[LoadQueue.scala 233:86:@38058.8]
  assign _T_92523 = _T_92522 | storeAddrNotKnownFlagsPReg_3_8; // @[LoadQueue.scala 233:86:@38059.8]
  assign _T_92524 = _T_92523 | storeAddrNotKnownFlagsPReg_3_9; // @[LoadQueue.scala 233:86:@38060.8]
  assign _T_92525 = _T_92524 | storeAddrNotKnownFlagsPReg_3_10; // @[LoadQueue.scala 233:86:@38061.8]
  assign _T_92526 = _T_92525 | storeAddrNotKnownFlagsPReg_3_11; // @[LoadQueue.scala 233:86:@38062.8]
  assign _T_92527 = _T_92526 | storeAddrNotKnownFlagsPReg_3_12; // @[LoadQueue.scala 233:86:@38063.8]
  assign _T_92528 = _T_92527 | storeAddrNotKnownFlagsPReg_3_13; // @[LoadQueue.scala 233:86:@38064.8]
  assign _T_92529 = _T_92528 | storeAddrNotKnownFlagsPReg_3_14; // @[LoadQueue.scala 233:86:@38065.8]
  assign _T_92530 = _T_92529 | storeAddrNotKnownFlagsPReg_3_15; // @[LoadQueue.scala 233:86:@38066.8]
  assign _T_92532 = _T_92530 == 1'h0; // @[LoadQueue.scala 233:38:@38067.8]
  assign _T_92551 = _T_88706 == 1'h0; // @[LoadQueue.scala 234:11:@38084.8]
  assign _T_92552 = _T_92532 & _T_92551; // @[LoadQueue.scala 233:103:@38085.8]
  assign _GEN_1980 = _T_92513 ? _T_92552 : 1'h0; // @[LoadQueue.scala 230:110:@38050.6]
  assign loadRequest_3 = _T_92505 ? _GEN_1980 : 1'h0; // @[LoadQueue.scala 229:71:@38044.4]
  assign _T_90468 = loadRequest_3 ? 16'h8 : _T_90467; // @[Mux.scala 31:69:@36533.4]
  assign _T_92420 = dataKnownPReg_2 == 1'h0; // @[LoadQueue.scala 229:41:@37960.4]
  assign _T_92421 = addrKnownPReg_2 & _T_92420; // @[LoadQueue.scala 229:38:@37961.4]
  assign _T_92423 = bypassInitiated_2 == 1'h0; // @[LoadQueue.scala 230:12:@37963.6]
  assign _T_92425 = prevPriorityRequest_2 == 1'h0; // @[LoadQueue.scala 230:46:@37964.6]
  assign _T_92426 = _T_92423 & _T_92425; // @[LoadQueue.scala 230:43:@37965.6]
  assign _T_92428 = dataKnown_2 == 1'h0; // @[LoadQueue.scala 230:84:@37966.6]
  assign _T_92429 = _T_92426 & _T_92428; // @[LoadQueue.scala 230:81:@37967.6]
  assign _T_92432 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[LoadQueue.scala 233:86:@37970.8]
  assign _T_92433 = _T_92432 | storeAddrNotKnownFlagsPReg_2_2; // @[LoadQueue.scala 233:86:@37971.8]
  assign _T_92434 = _T_92433 | storeAddrNotKnownFlagsPReg_2_3; // @[LoadQueue.scala 233:86:@37972.8]
  assign _T_92435 = _T_92434 | storeAddrNotKnownFlagsPReg_2_4; // @[LoadQueue.scala 233:86:@37973.8]
  assign _T_92436 = _T_92435 | storeAddrNotKnownFlagsPReg_2_5; // @[LoadQueue.scala 233:86:@37974.8]
  assign _T_92437 = _T_92436 | storeAddrNotKnownFlagsPReg_2_6; // @[LoadQueue.scala 233:86:@37975.8]
  assign _T_92438 = _T_92437 | storeAddrNotKnownFlagsPReg_2_7; // @[LoadQueue.scala 233:86:@37976.8]
  assign _T_92439 = _T_92438 | storeAddrNotKnownFlagsPReg_2_8; // @[LoadQueue.scala 233:86:@37977.8]
  assign _T_92440 = _T_92439 | storeAddrNotKnownFlagsPReg_2_9; // @[LoadQueue.scala 233:86:@37978.8]
  assign _T_92441 = _T_92440 | storeAddrNotKnownFlagsPReg_2_10; // @[LoadQueue.scala 233:86:@37979.8]
  assign _T_92442 = _T_92441 | storeAddrNotKnownFlagsPReg_2_11; // @[LoadQueue.scala 233:86:@37980.8]
  assign _T_92443 = _T_92442 | storeAddrNotKnownFlagsPReg_2_12; // @[LoadQueue.scala 233:86:@37981.8]
  assign _T_92444 = _T_92443 | storeAddrNotKnownFlagsPReg_2_13; // @[LoadQueue.scala 233:86:@37982.8]
  assign _T_92445 = _T_92444 | storeAddrNotKnownFlagsPReg_2_14; // @[LoadQueue.scala 233:86:@37983.8]
  assign _T_92446 = _T_92445 | storeAddrNotKnownFlagsPReg_2_15; // @[LoadQueue.scala 233:86:@37984.8]
  assign _T_92448 = _T_92446 == 1'h0; // @[LoadQueue.scala 233:38:@37985.8]
  assign _T_92467 = _T_88570 == 1'h0; // @[LoadQueue.scala 234:11:@38002.8]
  assign _T_92468 = _T_92448 & _T_92467; // @[LoadQueue.scala 233:103:@38003.8]
  assign _GEN_1976 = _T_92429 ? _T_92468 : 1'h0; // @[LoadQueue.scala 230:110:@37968.6]
  assign loadRequest_2 = _T_92421 ? _GEN_1976 : 1'h0; // @[LoadQueue.scala 229:71:@37962.4]
  assign _T_90469 = loadRequest_2 ? 16'h4 : _T_90468; // @[Mux.scala 31:69:@36534.4]
  assign _T_92336 = dataKnownPReg_1 == 1'h0; // @[LoadQueue.scala 229:41:@37878.4]
  assign _T_92337 = addrKnownPReg_1 & _T_92336; // @[LoadQueue.scala 229:38:@37879.4]
  assign _T_92339 = bypassInitiated_1 == 1'h0; // @[LoadQueue.scala 230:12:@37881.6]
  assign _T_92341 = prevPriorityRequest_1 == 1'h0; // @[LoadQueue.scala 230:46:@37882.6]
  assign _T_92342 = _T_92339 & _T_92341; // @[LoadQueue.scala 230:43:@37883.6]
  assign _T_92344 = dataKnown_1 == 1'h0; // @[LoadQueue.scala 230:84:@37884.6]
  assign _T_92345 = _T_92342 & _T_92344; // @[LoadQueue.scala 230:81:@37885.6]
  assign _T_92348 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[LoadQueue.scala 233:86:@37888.8]
  assign _T_92349 = _T_92348 | storeAddrNotKnownFlagsPReg_1_2; // @[LoadQueue.scala 233:86:@37889.8]
  assign _T_92350 = _T_92349 | storeAddrNotKnownFlagsPReg_1_3; // @[LoadQueue.scala 233:86:@37890.8]
  assign _T_92351 = _T_92350 | storeAddrNotKnownFlagsPReg_1_4; // @[LoadQueue.scala 233:86:@37891.8]
  assign _T_92352 = _T_92351 | storeAddrNotKnownFlagsPReg_1_5; // @[LoadQueue.scala 233:86:@37892.8]
  assign _T_92353 = _T_92352 | storeAddrNotKnownFlagsPReg_1_6; // @[LoadQueue.scala 233:86:@37893.8]
  assign _T_92354 = _T_92353 | storeAddrNotKnownFlagsPReg_1_7; // @[LoadQueue.scala 233:86:@37894.8]
  assign _T_92355 = _T_92354 | storeAddrNotKnownFlagsPReg_1_8; // @[LoadQueue.scala 233:86:@37895.8]
  assign _T_92356 = _T_92355 | storeAddrNotKnownFlagsPReg_1_9; // @[LoadQueue.scala 233:86:@37896.8]
  assign _T_92357 = _T_92356 | storeAddrNotKnownFlagsPReg_1_10; // @[LoadQueue.scala 233:86:@37897.8]
  assign _T_92358 = _T_92357 | storeAddrNotKnownFlagsPReg_1_11; // @[LoadQueue.scala 233:86:@37898.8]
  assign _T_92359 = _T_92358 | storeAddrNotKnownFlagsPReg_1_12; // @[LoadQueue.scala 233:86:@37899.8]
  assign _T_92360 = _T_92359 | storeAddrNotKnownFlagsPReg_1_13; // @[LoadQueue.scala 233:86:@37900.8]
  assign _T_92361 = _T_92360 | storeAddrNotKnownFlagsPReg_1_14; // @[LoadQueue.scala 233:86:@37901.8]
  assign _T_92362 = _T_92361 | storeAddrNotKnownFlagsPReg_1_15; // @[LoadQueue.scala 233:86:@37902.8]
  assign _T_92364 = _T_92362 == 1'h0; // @[LoadQueue.scala 233:38:@37903.8]
  assign _T_92383 = _T_88434 == 1'h0; // @[LoadQueue.scala 234:11:@37920.8]
  assign _T_92384 = _T_92364 & _T_92383; // @[LoadQueue.scala 233:103:@37921.8]
  assign _GEN_1972 = _T_92345 ? _T_92384 : 1'h0; // @[LoadQueue.scala 230:110:@37886.6]
  assign loadRequest_1 = _T_92337 ? _GEN_1972 : 1'h0; // @[LoadQueue.scala 229:71:@37880.4]
  assign _T_90470 = loadRequest_1 ? 16'h2 : _T_90469; // @[Mux.scala 31:69:@36535.4]
  assign _T_92252 = dataKnownPReg_0 == 1'h0; // @[LoadQueue.scala 229:41:@37796.4]
  assign _T_92253 = addrKnownPReg_0 & _T_92252; // @[LoadQueue.scala 229:38:@37797.4]
  assign _T_92255 = bypassInitiated_0 == 1'h0; // @[LoadQueue.scala 230:12:@37799.6]
  assign _T_92257 = prevPriorityRequest_0 == 1'h0; // @[LoadQueue.scala 230:46:@37800.6]
  assign _T_92258 = _T_92255 & _T_92257; // @[LoadQueue.scala 230:43:@37801.6]
  assign _T_92260 = dataKnown_0 == 1'h0; // @[LoadQueue.scala 230:84:@37802.6]
  assign _T_92261 = _T_92258 & _T_92260; // @[LoadQueue.scala 230:81:@37803.6]
  assign _T_92264 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[LoadQueue.scala 233:86:@37806.8]
  assign _T_92265 = _T_92264 | storeAddrNotKnownFlagsPReg_0_2; // @[LoadQueue.scala 233:86:@37807.8]
  assign _T_92266 = _T_92265 | storeAddrNotKnownFlagsPReg_0_3; // @[LoadQueue.scala 233:86:@37808.8]
  assign _T_92267 = _T_92266 | storeAddrNotKnownFlagsPReg_0_4; // @[LoadQueue.scala 233:86:@37809.8]
  assign _T_92268 = _T_92267 | storeAddrNotKnownFlagsPReg_0_5; // @[LoadQueue.scala 233:86:@37810.8]
  assign _T_92269 = _T_92268 | storeAddrNotKnownFlagsPReg_0_6; // @[LoadQueue.scala 233:86:@37811.8]
  assign _T_92270 = _T_92269 | storeAddrNotKnownFlagsPReg_0_7; // @[LoadQueue.scala 233:86:@37812.8]
  assign _T_92271 = _T_92270 | storeAddrNotKnownFlagsPReg_0_8; // @[LoadQueue.scala 233:86:@37813.8]
  assign _T_92272 = _T_92271 | storeAddrNotKnownFlagsPReg_0_9; // @[LoadQueue.scala 233:86:@37814.8]
  assign _T_92273 = _T_92272 | storeAddrNotKnownFlagsPReg_0_10; // @[LoadQueue.scala 233:86:@37815.8]
  assign _T_92274 = _T_92273 | storeAddrNotKnownFlagsPReg_0_11; // @[LoadQueue.scala 233:86:@37816.8]
  assign _T_92275 = _T_92274 | storeAddrNotKnownFlagsPReg_0_12; // @[LoadQueue.scala 233:86:@37817.8]
  assign _T_92276 = _T_92275 | storeAddrNotKnownFlagsPReg_0_13; // @[LoadQueue.scala 233:86:@37818.8]
  assign _T_92277 = _T_92276 | storeAddrNotKnownFlagsPReg_0_14; // @[LoadQueue.scala 233:86:@37819.8]
  assign _T_92278 = _T_92277 | storeAddrNotKnownFlagsPReg_0_15; // @[LoadQueue.scala 233:86:@37820.8]
  assign _T_92280 = _T_92278 == 1'h0; // @[LoadQueue.scala 233:38:@37821.8]
  assign _T_92299 = _T_88298 == 1'h0; // @[LoadQueue.scala 234:11:@37838.8]
  assign _T_92300 = _T_92280 & _T_92299; // @[LoadQueue.scala 233:103:@37839.8]
  assign _GEN_1968 = _T_92261 ? _T_92300 : 1'h0; // @[LoadQueue.scala 230:110:@37804.6]
  assign loadRequest_0 = _T_92253 ? _GEN_1968 : 1'h0; // @[LoadQueue.scala 229:71:@37798.4]
  assign _T_90471 = loadRequest_0 ? 16'h1 : _T_90470; // @[Mux.scala 31:69:@36536.4]
  assign _T_90472 = _T_90471[0]; // @[OneHot.scala 66:30:@36537.4]
  assign _T_90473 = _T_90471[1]; // @[OneHot.scala 66:30:@36538.4]
  assign _T_90474 = _T_90471[2]; // @[OneHot.scala 66:30:@36539.4]
  assign _T_90475 = _T_90471[3]; // @[OneHot.scala 66:30:@36540.4]
  assign _T_90476 = _T_90471[4]; // @[OneHot.scala 66:30:@36541.4]
  assign _T_90477 = _T_90471[5]; // @[OneHot.scala 66:30:@36542.4]
  assign _T_90478 = _T_90471[6]; // @[OneHot.scala 66:30:@36543.4]
  assign _T_90479 = _T_90471[7]; // @[OneHot.scala 66:30:@36544.4]
  assign _T_90480 = _T_90471[8]; // @[OneHot.scala 66:30:@36545.4]
  assign _T_90481 = _T_90471[9]; // @[OneHot.scala 66:30:@36546.4]
  assign _T_90482 = _T_90471[10]; // @[OneHot.scala 66:30:@36547.4]
  assign _T_90483 = _T_90471[11]; // @[OneHot.scala 66:30:@36548.4]
  assign _T_90484 = _T_90471[12]; // @[OneHot.scala 66:30:@36549.4]
  assign _T_90485 = _T_90471[13]; // @[OneHot.scala 66:30:@36550.4]
  assign _T_90486 = _T_90471[14]; // @[OneHot.scala 66:30:@36551.4]
  assign _T_90487 = _T_90471[15]; // @[OneHot.scala 66:30:@36552.4]
  assign _T_90528 = loadRequest_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36570.4]
  assign _T_90529 = loadRequest_15 ? 16'h4000 : _T_90528; // @[Mux.scala 31:69:@36571.4]
  assign _T_90530 = loadRequest_14 ? 16'h2000 : _T_90529; // @[Mux.scala 31:69:@36572.4]
  assign _T_90531 = loadRequest_13 ? 16'h1000 : _T_90530; // @[Mux.scala 31:69:@36573.4]
  assign _T_90532 = loadRequest_12 ? 16'h800 : _T_90531; // @[Mux.scala 31:69:@36574.4]
  assign _T_90533 = loadRequest_11 ? 16'h400 : _T_90532; // @[Mux.scala 31:69:@36575.4]
  assign _T_90534 = loadRequest_10 ? 16'h200 : _T_90533; // @[Mux.scala 31:69:@36576.4]
  assign _T_90535 = loadRequest_9 ? 16'h100 : _T_90534; // @[Mux.scala 31:69:@36577.4]
  assign _T_90536 = loadRequest_8 ? 16'h80 : _T_90535; // @[Mux.scala 31:69:@36578.4]
  assign _T_90537 = loadRequest_7 ? 16'h40 : _T_90536; // @[Mux.scala 31:69:@36579.4]
  assign _T_90538 = loadRequest_6 ? 16'h20 : _T_90537; // @[Mux.scala 31:69:@36580.4]
  assign _T_90539 = loadRequest_5 ? 16'h10 : _T_90538; // @[Mux.scala 31:69:@36581.4]
  assign _T_90540 = loadRequest_4 ? 16'h8 : _T_90539; // @[Mux.scala 31:69:@36582.4]
  assign _T_90541 = loadRequest_3 ? 16'h4 : _T_90540; // @[Mux.scala 31:69:@36583.4]
  assign _T_90542 = loadRequest_2 ? 16'h2 : _T_90541; // @[Mux.scala 31:69:@36584.4]
  assign _T_90543 = loadRequest_1 ? 16'h1 : _T_90542; // @[Mux.scala 31:69:@36585.4]
  assign _T_90544 = _T_90543[0]; // @[OneHot.scala 66:30:@36586.4]
  assign _T_90545 = _T_90543[1]; // @[OneHot.scala 66:30:@36587.4]
  assign _T_90546 = _T_90543[2]; // @[OneHot.scala 66:30:@36588.4]
  assign _T_90547 = _T_90543[3]; // @[OneHot.scala 66:30:@36589.4]
  assign _T_90548 = _T_90543[4]; // @[OneHot.scala 66:30:@36590.4]
  assign _T_90549 = _T_90543[5]; // @[OneHot.scala 66:30:@36591.4]
  assign _T_90550 = _T_90543[6]; // @[OneHot.scala 66:30:@36592.4]
  assign _T_90551 = _T_90543[7]; // @[OneHot.scala 66:30:@36593.4]
  assign _T_90552 = _T_90543[8]; // @[OneHot.scala 66:30:@36594.4]
  assign _T_90553 = _T_90543[9]; // @[OneHot.scala 66:30:@36595.4]
  assign _T_90554 = _T_90543[10]; // @[OneHot.scala 66:30:@36596.4]
  assign _T_90555 = _T_90543[11]; // @[OneHot.scala 66:30:@36597.4]
  assign _T_90556 = _T_90543[12]; // @[OneHot.scala 66:30:@36598.4]
  assign _T_90557 = _T_90543[13]; // @[OneHot.scala 66:30:@36599.4]
  assign _T_90558 = _T_90543[14]; // @[OneHot.scala 66:30:@36600.4]
  assign _T_90559 = _T_90543[15]; // @[OneHot.scala 66:30:@36601.4]
  assign _T_90600 = loadRequest_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36619.4]
  assign _T_90601 = loadRequest_0 ? 16'h4000 : _T_90600; // @[Mux.scala 31:69:@36620.4]
  assign _T_90602 = loadRequest_15 ? 16'h2000 : _T_90601; // @[Mux.scala 31:69:@36621.4]
  assign _T_90603 = loadRequest_14 ? 16'h1000 : _T_90602; // @[Mux.scala 31:69:@36622.4]
  assign _T_90604 = loadRequest_13 ? 16'h800 : _T_90603; // @[Mux.scala 31:69:@36623.4]
  assign _T_90605 = loadRequest_12 ? 16'h400 : _T_90604; // @[Mux.scala 31:69:@36624.4]
  assign _T_90606 = loadRequest_11 ? 16'h200 : _T_90605; // @[Mux.scala 31:69:@36625.4]
  assign _T_90607 = loadRequest_10 ? 16'h100 : _T_90606; // @[Mux.scala 31:69:@36626.4]
  assign _T_90608 = loadRequest_9 ? 16'h80 : _T_90607; // @[Mux.scala 31:69:@36627.4]
  assign _T_90609 = loadRequest_8 ? 16'h40 : _T_90608; // @[Mux.scala 31:69:@36628.4]
  assign _T_90610 = loadRequest_7 ? 16'h20 : _T_90609; // @[Mux.scala 31:69:@36629.4]
  assign _T_90611 = loadRequest_6 ? 16'h10 : _T_90610; // @[Mux.scala 31:69:@36630.4]
  assign _T_90612 = loadRequest_5 ? 16'h8 : _T_90611; // @[Mux.scala 31:69:@36631.4]
  assign _T_90613 = loadRequest_4 ? 16'h4 : _T_90612; // @[Mux.scala 31:69:@36632.4]
  assign _T_90614 = loadRequest_3 ? 16'h2 : _T_90613; // @[Mux.scala 31:69:@36633.4]
  assign _T_90615 = loadRequest_2 ? 16'h1 : _T_90614; // @[Mux.scala 31:69:@36634.4]
  assign _T_90616 = _T_90615[0]; // @[OneHot.scala 66:30:@36635.4]
  assign _T_90617 = _T_90615[1]; // @[OneHot.scala 66:30:@36636.4]
  assign _T_90618 = _T_90615[2]; // @[OneHot.scala 66:30:@36637.4]
  assign _T_90619 = _T_90615[3]; // @[OneHot.scala 66:30:@36638.4]
  assign _T_90620 = _T_90615[4]; // @[OneHot.scala 66:30:@36639.4]
  assign _T_90621 = _T_90615[5]; // @[OneHot.scala 66:30:@36640.4]
  assign _T_90622 = _T_90615[6]; // @[OneHot.scala 66:30:@36641.4]
  assign _T_90623 = _T_90615[7]; // @[OneHot.scala 66:30:@36642.4]
  assign _T_90624 = _T_90615[8]; // @[OneHot.scala 66:30:@36643.4]
  assign _T_90625 = _T_90615[9]; // @[OneHot.scala 66:30:@36644.4]
  assign _T_90626 = _T_90615[10]; // @[OneHot.scala 66:30:@36645.4]
  assign _T_90627 = _T_90615[11]; // @[OneHot.scala 66:30:@36646.4]
  assign _T_90628 = _T_90615[12]; // @[OneHot.scala 66:30:@36647.4]
  assign _T_90629 = _T_90615[13]; // @[OneHot.scala 66:30:@36648.4]
  assign _T_90630 = _T_90615[14]; // @[OneHot.scala 66:30:@36649.4]
  assign _T_90631 = _T_90615[15]; // @[OneHot.scala 66:30:@36650.4]
  assign _T_90672 = loadRequest_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36668.4]
  assign _T_90673 = loadRequest_1 ? 16'h4000 : _T_90672; // @[Mux.scala 31:69:@36669.4]
  assign _T_90674 = loadRequest_0 ? 16'h2000 : _T_90673; // @[Mux.scala 31:69:@36670.4]
  assign _T_90675 = loadRequest_15 ? 16'h1000 : _T_90674; // @[Mux.scala 31:69:@36671.4]
  assign _T_90676 = loadRequest_14 ? 16'h800 : _T_90675; // @[Mux.scala 31:69:@36672.4]
  assign _T_90677 = loadRequest_13 ? 16'h400 : _T_90676; // @[Mux.scala 31:69:@36673.4]
  assign _T_90678 = loadRequest_12 ? 16'h200 : _T_90677; // @[Mux.scala 31:69:@36674.4]
  assign _T_90679 = loadRequest_11 ? 16'h100 : _T_90678; // @[Mux.scala 31:69:@36675.4]
  assign _T_90680 = loadRequest_10 ? 16'h80 : _T_90679; // @[Mux.scala 31:69:@36676.4]
  assign _T_90681 = loadRequest_9 ? 16'h40 : _T_90680; // @[Mux.scala 31:69:@36677.4]
  assign _T_90682 = loadRequest_8 ? 16'h20 : _T_90681; // @[Mux.scala 31:69:@36678.4]
  assign _T_90683 = loadRequest_7 ? 16'h10 : _T_90682; // @[Mux.scala 31:69:@36679.4]
  assign _T_90684 = loadRequest_6 ? 16'h8 : _T_90683; // @[Mux.scala 31:69:@36680.4]
  assign _T_90685 = loadRequest_5 ? 16'h4 : _T_90684; // @[Mux.scala 31:69:@36681.4]
  assign _T_90686 = loadRequest_4 ? 16'h2 : _T_90685; // @[Mux.scala 31:69:@36682.4]
  assign _T_90687 = loadRequest_3 ? 16'h1 : _T_90686; // @[Mux.scala 31:69:@36683.4]
  assign _T_90688 = _T_90687[0]; // @[OneHot.scala 66:30:@36684.4]
  assign _T_90689 = _T_90687[1]; // @[OneHot.scala 66:30:@36685.4]
  assign _T_90690 = _T_90687[2]; // @[OneHot.scala 66:30:@36686.4]
  assign _T_90691 = _T_90687[3]; // @[OneHot.scala 66:30:@36687.4]
  assign _T_90692 = _T_90687[4]; // @[OneHot.scala 66:30:@36688.4]
  assign _T_90693 = _T_90687[5]; // @[OneHot.scala 66:30:@36689.4]
  assign _T_90694 = _T_90687[6]; // @[OneHot.scala 66:30:@36690.4]
  assign _T_90695 = _T_90687[7]; // @[OneHot.scala 66:30:@36691.4]
  assign _T_90696 = _T_90687[8]; // @[OneHot.scala 66:30:@36692.4]
  assign _T_90697 = _T_90687[9]; // @[OneHot.scala 66:30:@36693.4]
  assign _T_90698 = _T_90687[10]; // @[OneHot.scala 66:30:@36694.4]
  assign _T_90699 = _T_90687[11]; // @[OneHot.scala 66:30:@36695.4]
  assign _T_90700 = _T_90687[12]; // @[OneHot.scala 66:30:@36696.4]
  assign _T_90701 = _T_90687[13]; // @[OneHot.scala 66:30:@36697.4]
  assign _T_90702 = _T_90687[14]; // @[OneHot.scala 66:30:@36698.4]
  assign _T_90703 = _T_90687[15]; // @[OneHot.scala 66:30:@36699.4]
  assign _T_90744 = loadRequest_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36717.4]
  assign _T_90745 = loadRequest_2 ? 16'h4000 : _T_90744; // @[Mux.scala 31:69:@36718.4]
  assign _T_90746 = loadRequest_1 ? 16'h2000 : _T_90745; // @[Mux.scala 31:69:@36719.4]
  assign _T_90747 = loadRequest_0 ? 16'h1000 : _T_90746; // @[Mux.scala 31:69:@36720.4]
  assign _T_90748 = loadRequest_15 ? 16'h800 : _T_90747; // @[Mux.scala 31:69:@36721.4]
  assign _T_90749 = loadRequest_14 ? 16'h400 : _T_90748; // @[Mux.scala 31:69:@36722.4]
  assign _T_90750 = loadRequest_13 ? 16'h200 : _T_90749; // @[Mux.scala 31:69:@36723.4]
  assign _T_90751 = loadRequest_12 ? 16'h100 : _T_90750; // @[Mux.scala 31:69:@36724.4]
  assign _T_90752 = loadRequest_11 ? 16'h80 : _T_90751; // @[Mux.scala 31:69:@36725.4]
  assign _T_90753 = loadRequest_10 ? 16'h40 : _T_90752; // @[Mux.scala 31:69:@36726.4]
  assign _T_90754 = loadRequest_9 ? 16'h20 : _T_90753; // @[Mux.scala 31:69:@36727.4]
  assign _T_90755 = loadRequest_8 ? 16'h10 : _T_90754; // @[Mux.scala 31:69:@36728.4]
  assign _T_90756 = loadRequest_7 ? 16'h8 : _T_90755; // @[Mux.scala 31:69:@36729.4]
  assign _T_90757 = loadRequest_6 ? 16'h4 : _T_90756; // @[Mux.scala 31:69:@36730.4]
  assign _T_90758 = loadRequest_5 ? 16'h2 : _T_90757; // @[Mux.scala 31:69:@36731.4]
  assign _T_90759 = loadRequest_4 ? 16'h1 : _T_90758; // @[Mux.scala 31:69:@36732.4]
  assign _T_90760 = _T_90759[0]; // @[OneHot.scala 66:30:@36733.4]
  assign _T_90761 = _T_90759[1]; // @[OneHot.scala 66:30:@36734.4]
  assign _T_90762 = _T_90759[2]; // @[OneHot.scala 66:30:@36735.4]
  assign _T_90763 = _T_90759[3]; // @[OneHot.scala 66:30:@36736.4]
  assign _T_90764 = _T_90759[4]; // @[OneHot.scala 66:30:@36737.4]
  assign _T_90765 = _T_90759[5]; // @[OneHot.scala 66:30:@36738.4]
  assign _T_90766 = _T_90759[6]; // @[OneHot.scala 66:30:@36739.4]
  assign _T_90767 = _T_90759[7]; // @[OneHot.scala 66:30:@36740.4]
  assign _T_90768 = _T_90759[8]; // @[OneHot.scala 66:30:@36741.4]
  assign _T_90769 = _T_90759[9]; // @[OneHot.scala 66:30:@36742.4]
  assign _T_90770 = _T_90759[10]; // @[OneHot.scala 66:30:@36743.4]
  assign _T_90771 = _T_90759[11]; // @[OneHot.scala 66:30:@36744.4]
  assign _T_90772 = _T_90759[12]; // @[OneHot.scala 66:30:@36745.4]
  assign _T_90773 = _T_90759[13]; // @[OneHot.scala 66:30:@36746.4]
  assign _T_90774 = _T_90759[14]; // @[OneHot.scala 66:30:@36747.4]
  assign _T_90775 = _T_90759[15]; // @[OneHot.scala 66:30:@36748.4]
  assign _T_90816 = loadRequest_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36766.4]
  assign _T_90817 = loadRequest_3 ? 16'h4000 : _T_90816; // @[Mux.scala 31:69:@36767.4]
  assign _T_90818 = loadRequest_2 ? 16'h2000 : _T_90817; // @[Mux.scala 31:69:@36768.4]
  assign _T_90819 = loadRequest_1 ? 16'h1000 : _T_90818; // @[Mux.scala 31:69:@36769.4]
  assign _T_90820 = loadRequest_0 ? 16'h800 : _T_90819; // @[Mux.scala 31:69:@36770.4]
  assign _T_90821 = loadRequest_15 ? 16'h400 : _T_90820; // @[Mux.scala 31:69:@36771.4]
  assign _T_90822 = loadRequest_14 ? 16'h200 : _T_90821; // @[Mux.scala 31:69:@36772.4]
  assign _T_90823 = loadRequest_13 ? 16'h100 : _T_90822; // @[Mux.scala 31:69:@36773.4]
  assign _T_90824 = loadRequest_12 ? 16'h80 : _T_90823; // @[Mux.scala 31:69:@36774.4]
  assign _T_90825 = loadRequest_11 ? 16'h40 : _T_90824; // @[Mux.scala 31:69:@36775.4]
  assign _T_90826 = loadRequest_10 ? 16'h20 : _T_90825; // @[Mux.scala 31:69:@36776.4]
  assign _T_90827 = loadRequest_9 ? 16'h10 : _T_90826; // @[Mux.scala 31:69:@36777.4]
  assign _T_90828 = loadRequest_8 ? 16'h8 : _T_90827; // @[Mux.scala 31:69:@36778.4]
  assign _T_90829 = loadRequest_7 ? 16'h4 : _T_90828; // @[Mux.scala 31:69:@36779.4]
  assign _T_90830 = loadRequest_6 ? 16'h2 : _T_90829; // @[Mux.scala 31:69:@36780.4]
  assign _T_90831 = loadRequest_5 ? 16'h1 : _T_90830; // @[Mux.scala 31:69:@36781.4]
  assign _T_90832 = _T_90831[0]; // @[OneHot.scala 66:30:@36782.4]
  assign _T_90833 = _T_90831[1]; // @[OneHot.scala 66:30:@36783.4]
  assign _T_90834 = _T_90831[2]; // @[OneHot.scala 66:30:@36784.4]
  assign _T_90835 = _T_90831[3]; // @[OneHot.scala 66:30:@36785.4]
  assign _T_90836 = _T_90831[4]; // @[OneHot.scala 66:30:@36786.4]
  assign _T_90837 = _T_90831[5]; // @[OneHot.scala 66:30:@36787.4]
  assign _T_90838 = _T_90831[6]; // @[OneHot.scala 66:30:@36788.4]
  assign _T_90839 = _T_90831[7]; // @[OneHot.scala 66:30:@36789.4]
  assign _T_90840 = _T_90831[8]; // @[OneHot.scala 66:30:@36790.4]
  assign _T_90841 = _T_90831[9]; // @[OneHot.scala 66:30:@36791.4]
  assign _T_90842 = _T_90831[10]; // @[OneHot.scala 66:30:@36792.4]
  assign _T_90843 = _T_90831[11]; // @[OneHot.scala 66:30:@36793.4]
  assign _T_90844 = _T_90831[12]; // @[OneHot.scala 66:30:@36794.4]
  assign _T_90845 = _T_90831[13]; // @[OneHot.scala 66:30:@36795.4]
  assign _T_90846 = _T_90831[14]; // @[OneHot.scala 66:30:@36796.4]
  assign _T_90847 = _T_90831[15]; // @[OneHot.scala 66:30:@36797.4]
  assign _T_90888 = loadRequest_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36815.4]
  assign _T_90889 = loadRequest_4 ? 16'h4000 : _T_90888; // @[Mux.scala 31:69:@36816.4]
  assign _T_90890 = loadRequest_3 ? 16'h2000 : _T_90889; // @[Mux.scala 31:69:@36817.4]
  assign _T_90891 = loadRequest_2 ? 16'h1000 : _T_90890; // @[Mux.scala 31:69:@36818.4]
  assign _T_90892 = loadRequest_1 ? 16'h800 : _T_90891; // @[Mux.scala 31:69:@36819.4]
  assign _T_90893 = loadRequest_0 ? 16'h400 : _T_90892; // @[Mux.scala 31:69:@36820.4]
  assign _T_90894 = loadRequest_15 ? 16'h200 : _T_90893; // @[Mux.scala 31:69:@36821.4]
  assign _T_90895 = loadRequest_14 ? 16'h100 : _T_90894; // @[Mux.scala 31:69:@36822.4]
  assign _T_90896 = loadRequest_13 ? 16'h80 : _T_90895; // @[Mux.scala 31:69:@36823.4]
  assign _T_90897 = loadRequest_12 ? 16'h40 : _T_90896; // @[Mux.scala 31:69:@36824.4]
  assign _T_90898 = loadRequest_11 ? 16'h20 : _T_90897; // @[Mux.scala 31:69:@36825.4]
  assign _T_90899 = loadRequest_10 ? 16'h10 : _T_90898; // @[Mux.scala 31:69:@36826.4]
  assign _T_90900 = loadRequest_9 ? 16'h8 : _T_90899; // @[Mux.scala 31:69:@36827.4]
  assign _T_90901 = loadRequest_8 ? 16'h4 : _T_90900; // @[Mux.scala 31:69:@36828.4]
  assign _T_90902 = loadRequest_7 ? 16'h2 : _T_90901; // @[Mux.scala 31:69:@36829.4]
  assign _T_90903 = loadRequest_6 ? 16'h1 : _T_90902; // @[Mux.scala 31:69:@36830.4]
  assign _T_90904 = _T_90903[0]; // @[OneHot.scala 66:30:@36831.4]
  assign _T_90905 = _T_90903[1]; // @[OneHot.scala 66:30:@36832.4]
  assign _T_90906 = _T_90903[2]; // @[OneHot.scala 66:30:@36833.4]
  assign _T_90907 = _T_90903[3]; // @[OneHot.scala 66:30:@36834.4]
  assign _T_90908 = _T_90903[4]; // @[OneHot.scala 66:30:@36835.4]
  assign _T_90909 = _T_90903[5]; // @[OneHot.scala 66:30:@36836.4]
  assign _T_90910 = _T_90903[6]; // @[OneHot.scala 66:30:@36837.4]
  assign _T_90911 = _T_90903[7]; // @[OneHot.scala 66:30:@36838.4]
  assign _T_90912 = _T_90903[8]; // @[OneHot.scala 66:30:@36839.4]
  assign _T_90913 = _T_90903[9]; // @[OneHot.scala 66:30:@36840.4]
  assign _T_90914 = _T_90903[10]; // @[OneHot.scala 66:30:@36841.4]
  assign _T_90915 = _T_90903[11]; // @[OneHot.scala 66:30:@36842.4]
  assign _T_90916 = _T_90903[12]; // @[OneHot.scala 66:30:@36843.4]
  assign _T_90917 = _T_90903[13]; // @[OneHot.scala 66:30:@36844.4]
  assign _T_90918 = _T_90903[14]; // @[OneHot.scala 66:30:@36845.4]
  assign _T_90919 = _T_90903[15]; // @[OneHot.scala 66:30:@36846.4]
  assign _T_90960 = loadRequest_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36864.4]
  assign _T_90961 = loadRequest_5 ? 16'h4000 : _T_90960; // @[Mux.scala 31:69:@36865.4]
  assign _T_90962 = loadRequest_4 ? 16'h2000 : _T_90961; // @[Mux.scala 31:69:@36866.4]
  assign _T_90963 = loadRequest_3 ? 16'h1000 : _T_90962; // @[Mux.scala 31:69:@36867.4]
  assign _T_90964 = loadRequest_2 ? 16'h800 : _T_90963; // @[Mux.scala 31:69:@36868.4]
  assign _T_90965 = loadRequest_1 ? 16'h400 : _T_90964; // @[Mux.scala 31:69:@36869.4]
  assign _T_90966 = loadRequest_0 ? 16'h200 : _T_90965; // @[Mux.scala 31:69:@36870.4]
  assign _T_90967 = loadRequest_15 ? 16'h100 : _T_90966; // @[Mux.scala 31:69:@36871.4]
  assign _T_90968 = loadRequest_14 ? 16'h80 : _T_90967; // @[Mux.scala 31:69:@36872.4]
  assign _T_90969 = loadRequest_13 ? 16'h40 : _T_90968; // @[Mux.scala 31:69:@36873.4]
  assign _T_90970 = loadRequest_12 ? 16'h20 : _T_90969; // @[Mux.scala 31:69:@36874.4]
  assign _T_90971 = loadRequest_11 ? 16'h10 : _T_90970; // @[Mux.scala 31:69:@36875.4]
  assign _T_90972 = loadRequest_10 ? 16'h8 : _T_90971; // @[Mux.scala 31:69:@36876.4]
  assign _T_90973 = loadRequest_9 ? 16'h4 : _T_90972; // @[Mux.scala 31:69:@36877.4]
  assign _T_90974 = loadRequest_8 ? 16'h2 : _T_90973; // @[Mux.scala 31:69:@36878.4]
  assign _T_90975 = loadRequest_7 ? 16'h1 : _T_90974; // @[Mux.scala 31:69:@36879.4]
  assign _T_90976 = _T_90975[0]; // @[OneHot.scala 66:30:@36880.4]
  assign _T_90977 = _T_90975[1]; // @[OneHot.scala 66:30:@36881.4]
  assign _T_90978 = _T_90975[2]; // @[OneHot.scala 66:30:@36882.4]
  assign _T_90979 = _T_90975[3]; // @[OneHot.scala 66:30:@36883.4]
  assign _T_90980 = _T_90975[4]; // @[OneHot.scala 66:30:@36884.4]
  assign _T_90981 = _T_90975[5]; // @[OneHot.scala 66:30:@36885.4]
  assign _T_90982 = _T_90975[6]; // @[OneHot.scala 66:30:@36886.4]
  assign _T_90983 = _T_90975[7]; // @[OneHot.scala 66:30:@36887.4]
  assign _T_90984 = _T_90975[8]; // @[OneHot.scala 66:30:@36888.4]
  assign _T_90985 = _T_90975[9]; // @[OneHot.scala 66:30:@36889.4]
  assign _T_90986 = _T_90975[10]; // @[OneHot.scala 66:30:@36890.4]
  assign _T_90987 = _T_90975[11]; // @[OneHot.scala 66:30:@36891.4]
  assign _T_90988 = _T_90975[12]; // @[OneHot.scala 66:30:@36892.4]
  assign _T_90989 = _T_90975[13]; // @[OneHot.scala 66:30:@36893.4]
  assign _T_90990 = _T_90975[14]; // @[OneHot.scala 66:30:@36894.4]
  assign _T_90991 = _T_90975[15]; // @[OneHot.scala 66:30:@36895.4]
  assign _T_91032 = loadRequest_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36913.4]
  assign _T_91033 = loadRequest_6 ? 16'h4000 : _T_91032; // @[Mux.scala 31:69:@36914.4]
  assign _T_91034 = loadRequest_5 ? 16'h2000 : _T_91033; // @[Mux.scala 31:69:@36915.4]
  assign _T_91035 = loadRequest_4 ? 16'h1000 : _T_91034; // @[Mux.scala 31:69:@36916.4]
  assign _T_91036 = loadRequest_3 ? 16'h800 : _T_91035; // @[Mux.scala 31:69:@36917.4]
  assign _T_91037 = loadRequest_2 ? 16'h400 : _T_91036; // @[Mux.scala 31:69:@36918.4]
  assign _T_91038 = loadRequest_1 ? 16'h200 : _T_91037; // @[Mux.scala 31:69:@36919.4]
  assign _T_91039 = loadRequest_0 ? 16'h100 : _T_91038; // @[Mux.scala 31:69:@36920.4]
  assign _T_91040 = loadRequest_15 ? 16'h80 : _T_91039; // @[Mux.scala 31:69:@36921.4]
  assign _T_91041 = loadRequest_14 ? 16'h40 : _T_91040; // @[Mux.scala 31:69:@36922.4]
  assign _T_91042 = loadRequest_13 ? 16'h20 : _T_91041; // @[Mux.scala 31:69:@36923.4]
  assign _T_91043 = loadRequest_12 ? 16'h10 : _T_91042; // @[Mux.scala 31:69:@36924.4]
  assign _T_91044 = loadRequest_11 ? 16'h8 : _T_91043; // @[Mux.scala 31:69:@36925.4]
  assign _T_91045 = loadRequest_10 ? 16'h4 : _T_91044; // @[Mux.scala 31:69:@36926.4]
  assign _T_91046 = loadRequest_9 ? 16'h2 : _T_91045; // @[Mux.scala 31:69:@36927.4]
  assign _T_91047 = loadRequest_8 ? 16'h1 : _T_91046; // @[Mux.scala 31:69:@36928.4]
  assign _T_91048 = _T_91047[0]; // @[OneHot.scala 66:30:@36929.4]
  assign _T_91049 = _T_91047[1]; // @[OneHot.scala 66:30:@36930.4]
  assign _T_91050 = _T_91047[2]; // @[OneHot.scala 66:30:@36931.4]
  assign _T_91051 = _T_91047[3]; // @[OneHot.scala 66:30:@36932.4]
  assign _T_91052 = _T_91047[4]; // @[OneHot.scala 66:30:@36933.4]
  assign _T_91053 = _T_91047[5]; // @[OneHot.scala 66:30:@36934.4]
  assign _T_91054 = _T_91047[6]; // @[OneHot.scala 66:30:@36935.4]
  assign _T_91055 = _T_91047[7]; // @[OneHot.scala 66:30:@36936.4]
  assign _T_91056 = _T_91047[8]; // @[OneHot.scala 66:30:@36937.4]
  assign _T_91057 = _T_91047[9]; // @[OneHot.scala 66:30:@36938.4]
  assign _T_91058 = _T_91047[10]; // @[OneHot.scala 66:30:@36939.4]
  assign _T_91059 = _T_91047[11]; // @[OneHot.scala 66:30:@36940.4]
  assign _T_91060 = _T_91047[12]; // @[OneHot.scala 66:30:@36941.4]
  assign _T_91061 = _T_91047[13]; // @[OneHot.scala 66:30:@36942.4]
  assign _T_91062 = _T_91047[14]; // @[OneHot.scala 66:30:@36943.4]
  assign _T_91063 = _T_91047[15]; // @[OneHot.scala 66:30:@36944.4]
  assign _T_91104 = loadRequest_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36962.4]
  assign _T_91105 = loadRequest_7 ? 16'h4000 : _T_91104; // @[Mux.scala 31:69:@36963.4]
  assign _T_91106 = loadRequest_6 ? 16'h2000 : _T_91105; // @[Mux.scala 31:69:@36964.4]
  assign _T_91107 = loadRequest_5 ? 16'h1000 : _T_91106; // @[Mux.scala 31:69:@36965.4]
  assign _T_91108 = loadRequest_4 ? 16'h800 : _T_91107; // @[Mux.scala 31:69:@36966.4]
  assign _T_91109 = loadRequest_3 ? 16'h400 : _T_91108; // @[Mux.scala 31:69:@36967.4]
  assign _T_91110 = loadRequest_2 ? 16'h200 : _T_91109; // @[Mux.scala 31:69:@36968.4]
  assign _T_91111 = loadRequest_1 ? 16'h100 : _T_91110; // @[Mux.scala 31:69:@36969.4]
  assign _T_91112 = loadRequest_0 ? 16'h80 : _T_91111; // @[Mux.scala 31:69:@36970.4]
  assign _T_91113 = loadRequest_15 ? 16'h40 : _T_91112; // @[Mux.scala 31:69:@36971.4]
  assign _T_91114 = loadRequest_14 ? 16'h20 : _T_91113; // @[Mux.scala 31:69:@36972.4]
  assign _T_91115 = loadRequest_13 ? 16'h10 : _T_91114; // @[Mux.scala 31:69:@36973.4]
  assign _T_91116 = loadRequest_12 ? 16'h8 : _T_91115; // @[Mux.scala 31:69:@36974.4]
  assign _T_91117 = loadRequest_11 ? 16'h4 : _T_91116; // @[Mux.scala 31:69:@36975.4]
  assign _T_91118 = loadRequest_10 ? 16'h2 : _T_91117; // @[Mux.scala 31:69:@36976.4]
  assign _T_91119 = loadRequest_9 ? 16'h1 : _T_91118; // @[Mux.scala 31:69:@36977.4]
  assign _T_91120 = _T_91119[0]; // @[OneHot.scala 66:30:@36978.4]
  assign _T_91121 = _T_91119[1]; // @[OneHot.scala 66:30:@36979.4]
  assign _T_91122 = _T_91119[2]; // @[OneHot.scala 66:30:@36980.4]
  assign _T_91123 = _T_91119[3]; // @[OneHot.scala 66:30:@36981.4]
  assign _T_91124 = _T_91119[4]; // @[OneHot.scala 66:30:@36982.4]
  assign _T_91125 = _T_91119[5]; // @[OneHot.scala 66:30:@36983.4]
  assign _T_91126 = _T_91119[6]; // @[OneHot.scala 66:30:@36984.4]
  assign _T_91127 = _T_91119[7]; // @[OneHot.scala 66:30:@36985.4]
  assign _T_91128 = _T_91119[8]; // @[OneHot.scala 66:30:@36986.4]
  assign _T_91129 = _T_91119[9]; // @[OneHot.scala 66:30:@36987.4]
  assign _T_91130 = _T_91119[10]; // @[OneHot.scala 66:30:@36988.4]
  assign _T_91131 = _T_91119[11]; // @[OneHot.scala 66:30:@36989.4]
  assign _T_91132 = _T_91119[12]; // @[OneHot.scala 66:30:@36990.4]
  assign _T_91133 = _T_91119[13]; // @[OneHot.scala 66:30:@36991.4]
  assign _T_91134 = _T_91119[14]; // @[OneHot.scala 66:30:@36992.4]
  assign _T_91135 = _T_91119[15]; // @[OneHot.scala 66:30:@36993.4]
  assign _T_91176 = loadRequest_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37011.4]
  assign _T_91177 = loadRequest_8 ? 16'h4000 : _T_91176; // @[Mux.scala 31:69:@37012.4]
  assign _T_91178 = loadRequest_7 ? 16'h2000 : _T_91177; // @[Mux.scala 31:69:@37013.4]
  assign _T_91179 = loadRequest_6 ? 16'h1000 : _T_91178; // @[Mux.scala 31:69:@37014.4]
  assign _T_91180 = loadRequest_5 ? 16'h800 : _T_91179; // @[Mux.scala 31:69:@37015.4]
  assign _T_91181 = loadRequest_4 ? 16'h400 : _T_91180; // @[Mux.scala 31:69:@37016.4]
  assign _T_91182 = loadRequest_3 ? 16'h200 : _T_91181; // @[Mux.scala 31:69:@37017.4]
  assign _T_91183 = loadRequest_2 ? 16'h100 : _T_91182; // @[Mux.scala 31:69:@37018.4]
  assign _T_91184 = loadRequest_1 ? 16'h80 : _T_91183; // @[Mux.scala 31:69:@37019.4]
  assign _T_91185 = loadRequest_0 ? 16'h40 : _T_91184; // @[Mux.scala 31:69:@37020.4]
  assign _T_91186 = loadRequest_15 ? 16'h20 : _T_91185; // @[Mux.scala 31:69:@37021.4]
  assign _T_91187 = loadRequest_14 ? 16'h10 : _T_91186; // @[Mux.scala 31:69:@37022.4]
  assign _T_91188 = loadRequest_13 ? 16'h8 : _T_91187; // @[Mux.scala 31:69:@37023.4]
  assign _T_91189 = loadRequest_12 ? 16'h4 : _T_91188; // @[Mux.scala 31:69:@37024.4]
  assign _T_91190 = loadRequest_11 ? 16'h2 : _T_91189; // @[Mux.scala 31:69:@37025.4]
  assign _T_91191 = loadRequest_10 ? 16'h1 : _T_91190; // @[Mux.scala 31:69:@37026.4]
  assign _T_91192 = _T_91191[0]; // @[OneHot.scala 66:30:@37027.4]
  assign _T_91193 = _T_91191[1]; // @[OneHot.scala 66:30:@37028.4]
  assign _T_91194 = _T_91191[2]; // @[OneHot.scala 66:30:@37029.4]
  assign _T_91195 = _T_91191[3]; // @[OneHot.scala 66:30:@37030.4]
  assign _T_91196 = _T_91191[4]; // @[OneHot.scala 66:30:@37031.4]
  assign _T_91197 = _T_91191[5]; // @[OneHot.scala 66:30:@37032.4]
  assign _T_91198 = _T_91191[6]; // @[OneHot.scala 66:30:@37033.4]
  assign _T_91199 = _T_91191[7]; // @[OneHot.scala 66:30:@37034.4]
  assign _T_91200 = _T_91191[8]; // @[OneHot.scala 66:30:@37035.4]
  assign _T_91201 = _T_91191[9]; // @[OneHot.scala 66:30:@37036.4]
  assign _T_91202 = _T_91191[10]; // @[OneHot.scala 66:30:@37037.4]
  assign _T_91203 = _T_91191[11]; // @[OneHot.scala 66:30:@37038.4]
  assign _T_91204 = _T_91191[12]; // @[OneHot.scala 66:30:@37039.4]
  assign _T_91205 = _T_91191[13]; // @[OneHot.scala 66:30:@37040.4]
  assign _T_91206 = _T_91191[14]; // @[OneHot.scala 66:30:@37041.4]
  assign _T_91207 = _T_91191[15]; // @[OneHot.scala 66:30:@37042.4]
  assign _T_91248 = loadRequest_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37060.4]
  assign _T_91249 = loadRequest_9 ? 16'h4000 : _T_91248; // @[Mux.scala 31:69:@37061.4]
  assign _T_91250 = loadRequest_8 ? 16'h2000 : _T_91249; // @[Mux.scala 31:69:@37062.4]
  assign _T_91251 = loadRequest_7 ? 16'h1000 : _T_91250; // @[Mux.scala 31:69:@37063.4]
  assign _T_91252 = loadRequest_6 ? 16'h800 : _T_91251; // @[Mux.scala 31:69:@37064.4]
  assign _T_91253 = loadRequest_5 ? 16'h400 : _T_91252; // @[Mux.scala 31:69:@37065.4]
  assign _T_91254 = loadRequest_4 ? 16'h200 : _T_91253; // @[Mux.scala 31:69:@37066.4]
  assign _T_91255 = loadRequest_3 ? 16'h100 : _T_91254; // @[Mux.scala 31:69:@37067.4]
  assign _T_91256 = loadRequest_2 ? 16'h80 : _T_91255; // @[Mux.scala 31:69:@37068.4]
  assign _T_91257 = loadRequest_1 ? 16'h40 : _T_91256; // @[Mux.scala 31:69:@37069.4]
  assign _T_91258 = loadRequest_0 ? 16'h20 : _T_91257; // @[Mux.scala 31:69:@37070.4]
  assign _T_91259 = loadRequest_15 ? 16'h10 : _T_91258; // @[Mux.scala 31:69:@37071.4]
  assign _T_91260 = loadRequest_14 ? 16'h8 : _T_91259; // @[Mux.scala 31:69:@37072.4]
  assign _T_91261 = loadRequest_13 ? 16'h4 : _T_91260; // @[Mux.scala 31:69:@37073.4]
  assign _T_91262 = loadRequest_12 ? 16'h2 : _T_91261; // @[Mux.scala 31:69:@37074.4]
  assign _T_91263 = loadRequest_11 ? 16'h1 : _T_91262; // @[Mux.scala 31:69:@37075.4]
  assign _T_91264 = _T_91263[0]; // @[OneHot.scala 66:30:@37076.4]
  assign _T_91265 = _T_91263[1]; // @[OneHot.scala 66:30:@37077.4]
  assign _T_91266 = _T_91263[2]; // @[OneHot.scala 66:30:@37078.4]
  assign _T_91267 = _T_91263[3]; // @[OneHot.scala 66:30:@37079.4]
  assign _T_91268 = _T_91263[4]; // @[OneHot.scala 66:30:@37080.4]
  assign _T_91269 = _T_91263[5]; // @[OneHot.scala 66:30:@37081.4]
  assign _T_91270 = _T_91263[6]; // @[OneHot.scala 66:30:@37082.4]
  assign _T_91271 = _T_91263[7]; // @[OneHot.scala 66:30:@37083.4]
  assign _T_91272 = _T_91263[8]; // @[OneHot.scala 66:30:@37084.4]
  assign _T_91273 = _T_91263[9]; // @[OneHot.scala 66:30:@37085.4]
  assign _T_91274 = _T_91263[10]; // @[OneHot.scala 66:30:@37086.4]
  assign _T_91275 = _T_91263[11]; // @[OneHot.scala 66:30:@37087.4]
  assign _T_91276 = _T_91263[12]; // @[OneHot.scala 66:30:@37088.4]
  assign _T_91277 = _T_91263[13]; // @[OneHot.scala 66:30:@37089.4]
  assign _T_91278 = _T_91263[14]; // @[OneHot.scala 66:30:@37090.4]
  assign _T_91279 = _T_91263[15]; // @[OneHot.scala 66:30:@37091.4]
  assign _T_91320 = loadRequest_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37109.4]
  assign _T_91321 = loadRequest_10 ? 16'h4000 : _T_91320; // @[Mux.scala 31:69:@37110.4]
  assign _T_91322 = loadRequest_9 ? 16'h2000 : _T_91321; // @[Mux.scala 31:69:@37111.4]
  assign _T_91323 = loadRequest_8 ? 16'h1000 : _T_91322; // @[Mux.scala 31:69:@37112.4]
  assign _T_91324 = loadRequest_7 ? 16'h800 : _T_91323; // @[Mux.scala 31:69:@37113.4]
  assign _T_91325 = loadRequest_6 ? 16'h400 : _T_91324; // @[Mux.scala 31:69:@37114.4]
  assign _T_91326 = loadRequest_5 ? 16'h200 : _T_91325; // @[Mux.scala 31:69:@37115.4]
  assign _T_91327 = loadRequest_4 ? 16'h100 : _T_91326; // @[Mux.scala 31:69:@37116.4]
  assign _T_91328 = loadRequest_3 ? 16'h80 : _T_91327; // @[Mux.scala 31:69:@37117.4]
  assign _T_91329 = loadRequest_2 ? 16'h40 : _T_91328; // @[Mux.scala 31:69:@37118.4]
  assign _T_91330 = loadRequest_1 ? 16'h20 : _T_91329; // @[Mux.scala 31:69:@37119.4]
  assign _T_91331 = loadRequest_0 ? 16'h10 : _T_91330; // @[Mux.scala 31:69:@37120.4]
  assign _T_91332 = loadRequest_15 ? 16'h8 : _T_91331; // @[Mux.scala 31:69:@37121.4]
  assign _T_91333 = loadRequest_14 ? 16'h4 : _T_91332; // @[Mux.scala 31:69:@37122.4]
  assign _T_91334 = loadRequest_13 ? 16'h2 : _T_91333; // @[Mux.scala 31:69:@37123.4]
  assign _T_91335 = loadRequest_12 ? 16'h1 : _T_91334; // @[Mux.scala 31:69:@37124.4]
  assign _T_91336 = _T_91335[0]; // @[OneHot.scala 66:30:@37125.4]
  assign _T_91337 = _T_91335[1]; // @[OneHot.scala 66:30:@37126.4]
  assign _T_91338 = _T_91335[2]; // @[OneHot.scala 66:30:@37127.4]
  assign _T_91339 = _T_91335[3]; // @[OneHot.scala 66:30:@37128.4]
  assign _T_91340 = _T_91335[4]; // @[OneHot.scala 66:30:@37129.4]
  assign _T_91341 = _T_91335[5]; // @[OneHot.scala 66:30:@37130.4]
  assign _T_91342 = _T_91335[6]; // @[OneHot.scala 66:30:@37131.4]
  assign _T_91343 = _T_91335[7]; // @[OneHot.scala 66:30:@37132.4]
  assign _T_91344 = _T_91335[8]; // @[OneHot.scala 66:30:@37133.4]
  assign _T_91345 = _T_91335[9]; // @[OneHot.scala 66:30:@37134.4]
  assign _T_91346 = _T_91335[10]; // @[OneHot.scala 66:30:@37135.4]
  assign _T_91347 = _T_91335[11]; // @[OneHot.scala 66:30:@37136.4]
  assign _T_91348 = _T_91335[12]; // @[OneHot.scala 66:30:@37137.4]
  assign _T_91349 = _T_91335[13]; // @[OneHot.scala 66:30:@37138.4]
  assign _T_91350 = _T_91335[14]; // @[OneHot.scala 66:30:@37139.4]
  assign _T_91351 = _T_91335[15]; // @[OneHot.scala 66:30:@37140.4]
  assign _T_91392 = loadRequest_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37158.4]
  assign _T_91393 = loadRequest_11 ? 16'h4000 : _T_91392; // @[Mux.scala 31:69:@37159.4]
  assign _T_91394 = loadRequest_10 ? 16'h2000 : _T_91393; // @[Mux.scala 31:69:@37160.4]
  assign _T_91395 = loadRequest_9 ? 16'h1000 : _T_91394; // @[Mux.scala 31:69:@37161.4]
  assign _T_91396 = loadRequest_8 ? 16'h800 : _T_91395; // @[Mux.scala 31:69:@37162.4]
  assign _T_91397 = loadRequest_7 ? 16'h400 : _T_91396; // @[Mux.scala 31:69:@37163.4]
  assign _T_91398 = loadRequest_6 ? 16'h200 : _T_91397; // @[Mux.scala 31:69:@37164.4]
  assign _T_91399 = loadRequest_5 ? 16'h100 : _T_91398; // @[Mux.scala 31:69:@37165.4]
  assign _T_91400 = loadRequest_4 ? 16'h80 : _T_91399; // @[Mux.scala 31:69:@37166.4]
  assign _T_91401 = loadRequest_3 ? 16'h40 : _T_91400; // @[Mux.scala 31:69:@37167.4]
  assign _T_91402 = loadRequest_2 ? 16'h20 : _T_91401; // @[Mux.scala 31:69:@37168.4]
  assign _T_91403 = loadRequest_1 ? 16'h10 : _T_91402; // @[Mux.scala 31:69:@37169.4]
  assign _T_91404 = loadRequest_0 ? 16'h8 : _T_91403; // @[Mux.scala 31:69:@37170.4]
  assign _T_91405 = loadRequest_15 ? 16'h4 : _T_91404; // @[Mux.scala 31:69:@37171.4]
  assign _T_91406 = loadRequest_14 ? 16'h2 : _T_91405; // @[Mux.scala 31:69:@37172.4]
  assign _T_91407 = loadRequest_13 ? 16'h1 : _T_91406; // @[Mux.scala 31:69:@37173.4]
  assign _T_91408 = _T_91407[0]; // @[OneHot.scala 66:30:@37174.4]
  assign _T_91409 = _T_91407[1]; // @[OneHot.scala 66:30:@37175.4]
  assign _T_91410 = _T_91407[2]; // @[OneHot.scala 66:30:@37176.4]
  assign _T_91411 = _T_91407[3]; // @[OneHot.scala 66:30:@37177.4]
  assign _T_91412 = _T_91407[4]; // @[OneHot.scala 66:30:@37178.4]
  assign _T_91413 = _T_91407[5]; // @[OneHot.scala 66:30:@37179.4]
  assign _T_91414 = _T_91407[6]; // @[OneHot.scala 66:30:@37180.4]
  assign _T_91415 = _T_91407[7]; // @[OneHot.scala 66:30:@37181.4]
  assign _T_91416 = _T_91407[8]; // @[OneHot.scala 66:30:@37182.4]
  assign _T_91417 = _T_91407[9]; // @[OneHot.scala 66:30:@37183.4]
  assign _T_91418 = _T_91407[10]; // @[OneHot.scala 66:30:@37184.4]
  assign _T_91419 = _T_91407[11]; // @[OneHot.scala 66:30:@37185.4]
  assign _T_91420 = _T_91407[12]; // @[OneHot.scala 66:30:@37186.4]
  assign _T_91421 = _T_91407[13]; // @[OneHot.scala 66:30:@37187.4]
  assign _T_91422 = _T_91407[14]; // @[OneHot.scala 66:30:@37188.4]
  assign _T_91423 = _T_91407[15]; // @[OneHot.scala 66:30:@37189.4]
  assign _T_91464 = loadRequest_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37207.4]
  assign _T_91465 = loadRequest_12 ? 16'h4000 : _T_91464; // @[Mux.scala 31:69:@37208.4]
  assign _T_91466 = loadRequest_11 ? 16'h2000 : _T_91465; // @[Mux.scala 31:69:@37209.4]
  assign _T_91467 = loadRequest_10 ? 16'h1000 : _T_91466; // @[Mux.scala 31:69:@37210.4]
  assign _T_91468 = loadRequest_9 ? 16'h800 : _T_91467; // @[Mux.scala 31:69:@37211.4]
  assign _T_91469 = loadRequest_8 ? 16'h400 : _T_91468; // @[Mux.scala 31:69:@37212.4]
  assign _T_91470 = loadRequest_7 ? 16'h200 : _T_91469; // @[Mux.scala 31:69:@37213.4]
  assign _T_91471 = loadRequest_6 ? 16'h100 : _T_91470; // @[Mux.scala 31:69:@37214.4]
  assign _T_91472 = loadRequest_5 ? 16'h80 : _T_91471; // @[Mux.scala 31:69:@37215.4]
  assign _T_91473 = loadRequest_4 ? 16'h40 : _T_91472; // @[Mux.scala 31:69:@37216.4]
  assign _T_91474 = loadRequest_3 ? 16'h20 : _T_91473; // @[Mux.scala 31:69:@37217.4]
  assign _T_91475 = loadRequest_2 ? 16'h10 : _T_91474; // @[Mux.scala 31:69:@37218.4]
  assign _T_91476 = loadRequest_1 ? 16'h8 : _T_91475; // @[Mux.scala 31:69:@37219.4]
  assign _T_91477 = loadRequest_0 ? 16'h4 : _T_91476; // @[Mux.scala 31:69:@37220.4]
  assign _T_91478 = loadRequest_15 ? 16'h2 : _T_91477; // @[Mux.scala 31:69:@37221.4]
  assign _T_91479 = loadRequest_14 ? 16'h1 : _T_91478; // @[Mux.scala 31:69:@37222.4]
  assign _T_91480 = _T_91479[0]; // @[OneHot.scala 66:30:@37223.4]
  assign _T_91481 = _T_91479[1]; // @[OneHot.scala 66:30:@37224.4]
  assign _T_91482 = _T_91479[2]; // @[OneHot.scala 66:30:@37225.4]
  assign _T_91483 = _T_91479[3]; // @[OneHot.scala 66:30:@37226.4]
  assign _T_91484 = _T_91479[4]; // @[OneHot.scala 66:30:@37227.4]
  assign _T_91485 = _T_91479[5]; // @[OneHot.scala 66:30:@37228.4]
  assign _T_91486 = _T_91479[6]; // @[OneHot.scala 66:30:@37229.4]
  assign _T_91487 = _T_91479[7]; // @[OneHot.scala 66:30:@37230.4]
  assign _T_91488 = _T_91479[8]; // @[OneHot.scala 66:30:@37231.4]
  assign _T_91489 = _T_91479[9]; // @[OneHot.scala 66:30:@37232.4]
  assign _T_91490 = _T_91479[10]; // @[OneHot.scala 66:30:@37233.4]
  assign _T_91491 = _T_91479[11]; // @[OneHot.scala 66:30:@37234.4]
  assign _T_91492 = _T_91479[12]; // @[OneHot.scala 66:30:@37235.4]
  assign _T_91493 = _T_91479[13]; // @[OneHot.scala 66:30:@37236.4]
  assign _T_91494 = _T_91479[14]; // @[OneHot.scala 66:30:@37237.4]
  assign _T_91495 = _T_91479[15]; // @[OneHot.scala 66:30:@37238.4]
  assign _T_91536 = loadRequest_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37256.4]
  assign _T_91537 = loadRequest_13 ? 16'h4000 : _T_91536; // @[Mux.scala 31:69:@37257.4]
  assign _T_91538 = loadRequest_12 ? 16'h2000 : _T_91537; // @[Mux.scala 31:69:@37258.4]
  assign _T_91539 = loadRequest_11 ? 16'h1000 : _T_91538; // @[Mux.scala 31:69:@37259.4]
  assign _T_91540 = loadRequest_10 ? 16'h800 : _T_91539; // @[Mux.scala 31:69:@37260.4]
  assign _T_91541 = loadRequest_9 ? 16'h400 : _T_91540; // @[Mux.scala 31:69:@37261.4]
  assign _T_91542 = loadRequest_8 ? 16'h200 : _T_91541; // @[Mux.scala 31:69:@37262.4]
  assign _T_91543 = loadRequest_7 ? 16'h100 : _T_91542; // @[Mux.scala 31:69:@37263.4]
  assign _T_91544 = loadRequest_6 ? 16'h80 : _T_91543; // @[Mux.scala 31:69:@37264.4]
  assign _T_91545 = loadRequest_5 ? 16'h40 : _T_91544; // @[Mux.scala 31:69:@37265.4]
  assign _T_91546 = loadRequest_4 ? 16'h20 : _T_91545; // @[Mux.scala 31:69:@37266.4]
  assign _T_91547 = loadRequest_3 ? 16'h10 : _T_91546; // @[Mux.scala 31:69:@37267.4]
  assign _T_91548 = loadRequest_2 ? 16'h8 : _T_91547; // @[Mux.scala 31:69:@37268.4]
  assign _T_91549 = loadRequest_1 ? 16'h4 : _T_91548; // @[Mux.scala 31:69:@37269.4]
  assign _T_91550 = loadRequest_0 ? 16'h2 : _T_91549; // @[Mux.scala 31:69:@37270.4]
  assign _T_91551 = loadRequest_15 ? 16'h1 : _T_91550; // @[Mux.scala 31:69:@37271.4]
  assign _T_91552 = _T_91551[0]; // @[OneHot.scala 66:30:@37272.4]
  assign _T_91553 = _T_91551[1]; // @[OneHot.scala 66:30:@37273.4]
  assign _T_91554 = _T_91551[2]; // @[OneHot.scala 66:30:@37274.4]
  assign _T_91555 = _T_91551[3]; // @[OneHot.scala 66:30:@37275.4]
  assign _T_91556 = _T_91551[4]; // @[OneHot.scala 66:30:@37276.4]
  assign _T_91557 = _T_91551[5]; // @[OneHot.scala 66:30:@37277.4]
  assign _T_91558 = _T_91551[6]; // @[OneHot.scala 66:30:@37278.4]
  assign _T_91559 = _T_91551[7]; // @[OneHot.scala 66:30:@37279.4]
  assign _T_91560 = _T_91551[8]; // @[OneHot.scala 66:30:@37280.4]
  assign _T_91561 = _T_91551[9]; // @[OneHot.scala 66:30:@37281.4]
  assign _T_91562 = _T_91551[10]; // @[OneHot.scala 66:30:@37282.4]
  assign _T_91563 = _T_91551[11]; // @[OneHot.scala 66:30:@37283.4]
  assign _T_91564 = _T_91551[12]; // @[OneHot.scala 66:30:@37284.4]
  assign _T_91565 = _T_91551[13]; // @[OneHot.scala 66:30:@37285.4]
  assign _T_91566 = _T_91551[14]; // @[OneHot.scala 66:30:@37286.4]
  assign _T_91567 = _T_91551[15]; // @[OneHot.scala 66:30:@37287.4]
  assign _T_91632 = {_T_90479,_T_90478,_T_90477,_T_90476,_T_90475,_T_90474,_T_90473,_T_90472}; // @[Mux.scala 19:72:@37311.4]
  assign _T_91640 = {_T_90487,_T_90486,_T_90485,_T_90484,_T_90483,_T_90482,_T_90481,_T_90480,_T_91632}; // @[Mux.scala 19:72:@37319.4]
  assign _T_91642 = _T_90400 ? _T_91640 : 16'h0; // @[Mux.scala 19:72:@37320.4]
  assign _T_91649 = {_T_90550,_T_90549,_T_90548,_T_90547,_T_90546,_T_90545,_T_90544,_T_90559}; // @[Mux.scala 19:72:@37327.4]
  assign _T_91657 = {_T_90558,_T_90557,_T_90556,_T_90555,_T_90554,_T_90553,_T_90552,_T_90551,_T_91649}; // @[Mux.scala 19:72:@37335.4]
  assign _T_91659 = _T_90401 ? _T_91657 : 16'h0; // @[Mux.scala 19:72:@37336.4]
  assign _T_91666 = {_T_90621,_T_90620,_T_90619,_T_90618,_T_90617,_T_90616,_T_90631,_T_90630}; // @[Mux.scala 19:72:@37343.4]
  assign _T_91674 = {_T_90629,_T_90628,_T_90627,_T_90626,_T_90625,_T_90624,_T_90623,_T_90622,_T_91666}; // @[Mux.scala 19:72:@37351.4]
  assign _T_91676 = _T_90402 ? _T_91674 : 16'h0; // @[Mux.scala 19:72:@37352.4]
  assign _T_91683 = {_T_90692,_T_90691,_T_90690,_T_90689,_T_90688,_T_90703,_T_90702,_T_90701}; // @[Mux.scala 19:72:@37359.4]
  assign _T_91691 = {_T_90700,_T_90699,_T_90698,_T_90697,_T_90696,_T_90695,_T_90694,_T_90693,_T_91683}; // @[Mux.scala 19:72:@37367.4]
  assign _T_91693 = _T_90403 ? _T_91691 : 16'h0; // @[Mux.scala 19:72:@37368.4]
  assign _T_91700 = {_T_90763,_T_90762,_T_90761,_T_90760,_T_90775,_T_90774,_T_90773,_T_90772}; // @[Mux.scala 19:72:@37375.4]
  assign _T_91708 = {_T_90771,_T_90770,_T_90769,_T_90768,_T_90767,_T_90766,_T_90765,_T_90764,_T_91700}; // @[Mux.scala 19:72:@37383.4]
  assign _T_91710 = _T_90404 ? _T_91708 : 16'h0; // @[Mux.scala 19:72:@37384.4]
  assign _T_91717 = {_T_90834,_T_90833,_T_90832,_T_90847,_T_90846,_T_90845,_T_90844,_T_90843}; // @[Mux.scala 19:72:@37391.4]
  assign _T_91725 = {_T_90842,_T_90841,_T_90840,_T_90839,_T_90838,_T_90837,_T_90836,_T_90835,_T_91717}; // @[Mux.scala 19:72:@37399.4]
  assign _T_91727 = _T_90405 ? _T_91725 : 16'h0; // @[Mux.scala 19:72:@37400.4]
  assign _T_91734 = {_T_90905,_T_90904,_T_90919,_T_90918,_T_90917,_T_90916,_T_90915,_T_90914}; // @[Mux.scala 19:72:@37407.4]
  assign _T_91742 = {_T_90913,_T_90912,_T_90911,_T_90910,_T_90909,_T_90908,_T_90907,_T_90906,_T_91734}; // @[Mux.scala 19:72:@37415.4]
  assign _T_91744 = _T_90406 ? _T_91742 : 16'h0; // @[Mux.scala 19:72:@37416.4]
  assign _T_91751 = {_T_90976,_T_90991,_T_90990,_T_90989,_T_90988,_T_90987,_T_90986,_T_90985}; // @[Mux.scala 19:72:@37423.4]
  assign _T_91759 = {_T_90984,_T_90983,_T_90982,_T_90981,_T_90980,_T_90979,_T_90978,_T_90977,_T_91751}; // @[Mux.scala 19:72:@37431.4]
  assign _T_91761 = _T_90407 ? _T_91759 : 16'h0; // @[Mux.scala 19:72:@37432.4]
  assign _T_91768 = {_T_91063,_T_91062,_T_91061,_T_91060,_T_91059,_T_91058,_T_91057,_T_91056}; // @[Mux.scala 19:72:@37439.4]
  assign _T_91776 = {_T_91055,_T_91054,_T_91053,_T_91052,_T_91051,_T_91050,_T_91049,_T_91048,_T_91768}; // @[Mux.scala 19:72:@37447.4]
  assign _T_91778 = _T_90408 ? _T_91776 : 16'h0; // @[Mux.scala 19:72:@37448.4]
  assign _T_91785 = {_T_91134,_T_91133,_T_91132,_T_91131,_T_91130,_T_91129,_T_91128,_T_91127}; // @[Mux.scala 19:72:@37455.4]
  assign _T_91793 = {_T_91126,_T_91125,_T_91124,_T_91123,_T_91122,_T_91121,_T_91120,_T_91135,_T_91785}; // @[Mux.scala 19:72:@37463.4]
  assign _T_91795 = _T_90409 ? _T_91793 : 16'h0; // @[Mux.scala 19:72:@37464.4]
  assign _T_91802 = {_T_91205,_T_91204,_T_91203,_T_91202,_T_91201,_T_91200,_T_91199,_T_91198}; // @[Mux.scala 19:72:@37471.4]
  assign _T_91810 = {_T_91197,_T_91196,_T_91195,_T_91194,_T_91193,_T_91192,_T_91207,_T_91206,_T_91802}; // @[Mux.scala 19:72:@37479.4]
  assign _T_91812 = _T_90410 ? _T_91810 : 16'h0; // @[Mux.scala 19:72:@37480.4]
  assign _T_91819 = {_T_91276,_T_91275,_T_91274,_T_91273,_T_91272,_T_91271,_T_91270,_T_91269}; // @[Mux.scala 19:72:@37487.4]
  assign _T_91827 = {_T_91268,_T_91267,_T_91266,_T_91265,_T_91264,_T_91279,_T_91278,_T_91277,_T_91819}; // @[Mux.scala 19:72:@37495.4]
  assign _T_91829 = _T_90411 ? _T_91827 : 16'h0; // @[Mux.scala 19:72:@37496.4]
  assign _T_91836 = {_T_91347,_T_91346,_T_91345,_T_91344,_T_91343,_T_91342,_T_91341,_T_91340}; // @[Mux.scala 19:72:@37503.4]
  assign _T_91844 = {_T_91339,_T_91338,_T_91337,_T_91336,_T_91351,_T_91350,_T_91349,_T_91348,_T_91836}; // @[Mux.scala 19:72:@37511.4]
  assign _T_91846 = _T_90412 ? _T_91844 : 16'h0; // @[Mux.scala 19:72:@37512.4]
  assign _T_91853 = {_T_91418,_T_91417,_T_91416,_T_91415,_T_91414,_T_91413,_T_91412,_T_91411}; // @[Mux.scala 19:72:@37519.4]
  assign _T_91861 = {_T_91410,_T_91409,_T_91408,_T_91423,_T_91422,_T_91421,_T_91420,_T_91419,_T_91853}; // @[Mux.scala 19:72:@37527.4]
  assign _T_91863 = _T_90413 ? _T_91861 : 16'h0; // @[Mux.scala 19:72:@37528.4]
  assign _T_91870 = {_T_91489,_T_91488,_T_91487,_T_91486,_T_91485,_T_91484,_T_91483,_T_91482}; // @[Mux.scala 19:72:@37535.4]
  assign _T_91878 = {_T_91481,_T_91480,_T_91495,_T_91494,_T_91493,_T_91492,_T_91491,_T_91490,_T_91870}; // @[Mux.scala 19:72:@37543.4]
  assign _T_91880 = _T_90414 ? _T_91878 : 16'h0; // @[Mux.scala 19:72:@37544.4]
  assign _T_91887 = {_T_91560,_T_91559,_T_91558,_T_91557,_T_91556,_T_91555,_T_91554,_T_91553}; // @[Mux.scala 19:72:@37551.4]
  assign _T_91895 = {_T_91552,_T_91567,_T_91566,_T_91565,_T_91564,_T_91563,_T_91562,_T_91561,_T_91887}; // @[Mux.scala 19:72:@37559.4]
  assign _T_91897 = _T_90415 ? _T_91895 : 16'h0; // @[Mux.scala 19:72:@37560.4]
  assign _T_91898 = _T_91642 | _T_91659; // @[Mux.scala 19:72:@37561.4]
  assign _T_91899 = _T_91898 | _T_91676; // @[Mux.scala 19:72:@37562.4]
  assign _T_91900 = _T_91899 | _T_91693; // @[Mux.scala 19:72:@37563.4]
  assign _T_91901 = _T_91900 | _T_91710; // @[Mux.scala 19:72:@37564.4]
  assign _T_91902 = _T_91901 | _T_91727; // @[Mux.scala 19:72:@37565.4]
  assign _T_91903 = _T_91902 | _T_91744; // @[Mux.scala 19:72:@37566.4]
  assign _T_91904 = _T_91903 | _T_91761; // @[Mux.scala 19:72:@37567.4]
  assign _T_91905 = _T_91904 | _T_91778; // @[Mux.scala 19:72:@37568.4]
  assign _T_91906 = _T_91905 | _T_91795; // @[Mux.scala 19:72:@37569.4]
  assign _T_91907 = _T_91906 | _T_91812; // @[Mux.scala 19:72:@37570.4]
  assign _T_91908 = _T_91907 | _T_91829; // @[Mux.scala 19:72:@37571.4]
  assign _T_91909 = _T_91908 | _T_91846; // @[Mux.scala 19:72:@37572.4]
  assign _T_91910 = _T_91909 | _T_91863; // @[Mux.scala 19:72:@37573.4]
  assign _T_91911 = _T_91910 | _T_91880; // @[Mux.scala 19:72:@37574.4]
  assign _T_91912 = _T_91911 | _T_91897; // @[Mux.scala 19:72:@37575.4]
  assign priorityLoadRequest_0 = _T_91912[0]; // @[Mux.scala 19:72:@37579.4]
  assign priorityLoadRequest_1 = _T_91912[1]; // @[Mux.scala 19:72:@37581.4]
  assign priorityLoadRequest_2 = _T_91912[2]; // @[Mux.scala 19:72:@37583.4]
  assign priorityLoadRequest_3 = _T_91912[3]; // @[Mux.scala 19:72:@37585.4]
  assign priorityLoadRequest_4 = _T_91912[4]; // @[Mux.scala 19:72:@37587.4]
  assign priorityLoadRequest_5 = _T_91912[5]; // @[Mux.scala 19:72:@37589.4]
  assign priorityLoadRequest_6 = _T_91912[6]; // @[Mux.scala 19:72:@37591.4]
  assign priorityLoadRequest_7 = _T_91912[7]; // @[Mux.scala 19:72:@37593.4]
  assign priorityLoadRequest_8 = _T_91912[8]; // @[Mux.scala 19:72:@37595.4]
  assign priorityLoadRequest_9 = _T_91912[9]; // @[Mux.scala 19:72:@37597.4]
  assign priorityLoadRequest_10 = _T_91912[10]; // @[Mux.scala 19:72:@37599.4]
  assign priorityLoadRequest_11 = _T_91912[11]; // @[Mux.scala 19:72:@37601.4]
  assign priorityLoadRequest_12 = _T_91912[12]; // @[Mux.scala 19:72:@37603.4]
  assign priorityLoadRequest_13 = _T_91912[13]; // @[Mux.scala 19:72:@37605.4]
  assign priorityLoadRequest_14 = _T_91912[14]; // @[Mux.scala 19:72:@37607.4]
  assign priorityLoadRequest_15 = _T_91912[15]; // @[Mux.scala 19:72:@37609.4]
  assign _GEN_1920 = io_memIsReadyForLoads ? priorityLoadRequest_0 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1921 = io_memIsReadyForLoads ? priorityLoadRequest_1 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1922 = io_memIsReadyForLoads ? priorityLoadRequest_2 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1923 = io_memIsReadyForLoads ? priorityLoadRequest_3 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1924 = io_memIsReadyForLoads ? priorityLoadRequest_4 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1925 = io_memIsReadyForLoads ? priorityLoadRequest_5 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1926 = io_memIsReadyForLoads ? priorityLoadRequest_6 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1927 = io_memIsReadyForLoads ? priorityLoadRequest_7 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1928 = io_memIsReadyForLoads ? priorityLoadRequest_8 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1929 = io_memIsReadyForLoads ? priorityLoadRequest_9 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1930 = io_memIsReadyForLoads ? priorityLoadRequest_10 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1931 = io_memIsReadyForLoads ? priorityLoadRequest_11 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1932 = io_memIsReadyForLoads ? priorityLoadRequest_12 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1933 = io_memIsReadyForLoads ? priorityLoadRequest_13 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1934 = io_memIsReadyForLoads ? priorityLoadRequest_14 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _GEN_1935 = io_memIsReadyForLoads ? priorityLoadRequest_15 : 1'h0; // @[LoadQueue.scala 208:31:@37629.4]
  assign _T_92307 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[LoadQueue.scala 238:58:@37847.8]
  assign _T_92315 = {storeAddrNotKnownFlagsPReg_0_15,storeAddrNotKnownFlagsPReg_0_14,storeAddrNotKnownFlagsPReg_0_13,storeAddrNotKnownFlagsPReg_0_12,storeAddrNotKnownFlagsPReg_0_11,storeAddrNotKnownFlagsPReg_0_10,storeAddrNotKnownFlagsPReg_0_9,storeAddrNotKnownFlagsPReg_0_8,_T_92307}; // @[LoadQueue.scala 238:58:@37855.8]
  assign _T_92322 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[LoadQueue.scala 238:96:@37862.8]
  assign _T_92330 = {lastConflict_0_15,lastConflict_0_14,lastConflict_0_13,lastConflict_0_12,lastConflict_0_11,lastConflict_0_10,lastConflict_0_9,lastConflict_0_8,_T_92322}; // @[LoadQueue.scala 238:96:@37870.8]
  assign _T_92331 = _T_92315 < _T_92330; // @[LoadQueue.scala 238:61:@37871.8]
  assign _T_92332 = canBypass_0 & _T_92331; // @[LoadQueue.scala 237:64:@37872.8]
  assign _GEN_1969 = _T_92261 ? _T_92332 : 1'h0; // @[LoadQueue.scala 230:110:@37804.6]
  assign bypassRequest_0 = _T_92253 ? _GEN_1969 : 1'h0; // @[LoadQueue.scala 229:71:@37798.4]
  assign _GEN_1936 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[LoadQueue.scala 217:34:@37686.6]
  assign _GEN_1937 = initBits_0 ? 1'h0 : _GEN_1936; // @[LoadQueue.scala 215:23:@37682.4]
  assign _T_92391 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[LoadQueue.scala 238:58:@37929.8]
  assign _T_92399 = {storeAddrNotKnownFlagsPReg_1_15,storeAddrNotKnownFlagsPReg_1_14,storeAddrNotKnownFlagsPReg_1_13,storeAddrNotKnownFlagsPReg_1_12,storeAddrNotKnownFlagsPReg_1_11,storeAddrNotKnownFlagsPReg_1_10,storeAddrNotKnownFlagsPReg_1_9,storeAddrNotKnownFlagsPReg_1_8,_T_92391}; // @[LoadQueue.scala 238:58:@37937.8]
  assign _T_92406 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[LoadQueue.scala 238:96:@37944.8]
  assign _T_92414 = {lastConflict_1_15,lastConflict_1_14,lastConflict_1_13,lastConflict_1_12,lastConflict_1_11,lastConflict_1_10,lastConflict_1_9,lastConflict_1_8,_T_92406}; // @[LoadQueue.scala 238:96:@37952.8]
  assign _T_92415 = _T_92399 < _T_92414; // @[LoadQueue.scala 238:61:@37953.8]
  assign _T_92416 = canBypass_1 & _T_92415; // @[LoadQueue.scala 237:64:@37954.8]
  assign _GEN_1973 = _T_92345 ? _T_92416 : 1'h0; // @[LoadQueue.scala 230:110:@37886.6]
  assign bypassRequest_1 = _T_92337 ? _GEN_1973 : 1'h0; // @[LoadQueue.scala 229:71:@37880.4]
  assign _GEN_1938 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[LoadQueue.scala 217:34:@37693.6]
  assign _GEN_1939 = initBits_1 ? 1'h0 : _GEN_1938; // @[LoadQueue.scala 215:23:@37689.4]
  assign _T_92475 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[LoadQueue.scala 238:58:@38011.8]
  assign _T_92483 = {storeAddrNotKnownFlagsPReg_2_15,storeAddrNotKnownFlagsPReg_2_14,storeAddrNotKnownFlagsPReg_2_13,storeAddrNotKnownFlagsPReg_2_12,storeAddrNotKnownFlagsPReg_2_11,storeAddrNotKnownFlagsPReg_2_10,storeAddrNotKnownFlagsPReg_2_9,storeAddrNotKnownFlagsPReg_2_8,_T_92475}; // @[LoadQueue.scala 238:58:@38019.8]
  assign _T_92490 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[LoadQueue.scala 238:96:@38026.8]
  assign _T_92498 = {lastConflict_2_15,lastConflict_2_14,lastConflict_2_13,lastConflict_2_12,lastConflict_2_11,lastConflict_2_10,lastConflict_2_9,lastConflict_2_8,_T_92490}; // @[LoadQueue.scala 238:96:@38034.8]
  assign _T_92499 = _T_92483 < _T_92498; // @[LoadQueue.scala 238:61:@38035.8]
  assign _T_92500 = canBypass_2 & _T_92499; // @[LoadQueue.scala 237:64:@38036.8]
  assign _GEN_1977 = _T_92429 ? _T_92500 : 1'h0; // @[LoadQueue.scala 230:110:@37968.6]
  assign bypassRequest_2 = _T_92421 ? _GEN_1977 : 1'h0; // @[LoadQueue.scala 229:71:@37962.4]
  assign _GEN_1940 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[LoadQueue.scala 217:34:@37700.6]
  assign _GEN_1941 = initBits_2 ? 1'h0 : _GEN_1940; // @[LoadQueue.scala 215:23:@37696.4]
  assign _T_92559 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[LoadQueue.scala 238:58:@38093.8]
  assign _T_92567 = {storeAddrNotKnownFlagsPReg_3_15,storeAddrNotKnownFlagsPReg_3_14,storeAddrNotKnownFlagsPReg_3_13,storeAddrNotKnownFlagsPReg_3_12,storeAddrNotKnownFlagsPReg_3_11,storeAddrNotKnownFlagsPReg_3_10,storeAddrNotKnownFlagsPReg_3_9,storeAddrNotKnownFlagsPReg_3_8,_T_92559}; // @[LoadQueue.scala 238:58:@38101.8]
  assign _T_92574 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[LoadQueue.scala 238:96:@38108.8]
  assign _T_92582 = {lastConflict_3_15,lastConflict_3_14,lastConflict_3_13,lastConflict_3_12,lastConflict_3_11,lastConflict_3_10,lastConflict_3_9,lastConflict_3_8,_T_92574}; // @[LoadQueue.scala 238:96:@38116.8]
  assign _T_92583 = _T_92567 < _T_92582; // @[LoadQueue.scala 238:61:@38117.8]
  assign _T_92584 = canBypass_3 & _T_92583; // @[LoadQueue.scala 237:64:@38118.8]
  assign _GEN_1981 = _T_92513 ? _T_92584 : 1'h0; // @[LoadQueue.scala 230:110:@38050.6]
  assign bypassRequest_3 = _T_92505 ? _GEN_1981 : 1'h0; // @[LoadQueue.scala 229:71:@38044.4]
  assign _GEN_1942 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[LoadQueue.scala 217:34:@37707.6]
  assign _GEN_1943 = initBits_3 ? 1'h0 : _GEN_1942; // @[LoadQueue.scala 215:23:@37703.4]
  assign _T_92643 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[LoadQueue.scala 238:58:@38175.8]
  assign _T_92651 = {storeAddrNotKnownFlagsPReg_4_15,storeAddrNotKnownFlagsPReg_4_14,storeAddrNotKnownFlagsPReg_4_13,storeAddrNotKnownFlagsPReg_4_12,storeAddrNotKnownFlagsPReg_4_11,storeAddrNotKnownFlagsPReg_4_10,storeAddrNotKnownFlagsPReg_4_9,storeAddrNotKnownFlagsPReg_4_8,_T_92643}; // @[LoadQueue.scala 238:58:@38183.8]
  assign _T_92658 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[LoadQueue.scala 238:96:@38190.8]
  assign _T_92666 = {lastConflict_4_15,lastConflict_4_14,lastConflict_4_13,lastConflict_4_12,lastConflict_4_11,lastConflict_4_10,lastConflict_4_9,lastConflict_4_8,_T_92658}; // @[LoadQueue.scala 238:96:@38198.8]
  assign _T_92667 = _T_92651 < _T_92666; // @[LoadQueue.scala 238:61:@38199.8]
  assign _T_92668 = canBypass_4 & _T_92667; // @[LoadQueue.scala 237:64:@38200.8]
  assign _GEN_1985 = _T_92597 ? _T_92668 : 1'h0; // @[LoadQueue.scala 230:110:@38132.6]
  assign bypassRequest_4 = _T_92589 ? _GEN_1985 : 1'h0; // @[LoadQueue.scala 229:71:@38126.4]
  assign _GEN_1944 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[LoadQueue.scala 217:34:@37714.6]
  assign _GEN_1945 = initBits_4 ? 1'h0 : _GEN_1944; // @[LoadQueue.scala 215:23:@37710.4]
  assign _T_92727 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[LoadQueue.scala 238:58:@38257.8]
  assign _T_92735 = {storeAddrNotKnownFlagsPReg_5_15,storeAddrNotKnownFlagsPReg_5_14,storeAddrNotKnownFlagsPReg_5_13,storeAddrNotKnownFlagsPReg_5_12,storeAddrNotKnownFlagsPReg_5_11,storeAddrNotKnownFlagsPReg_5_10,storeAddrNotKnownFlagsPReg_5_9,storeAddrNotKnownFlagsPReg_5_8,_T_92727}; // @[LoadQueue.scala 238:58:@38265.8]
  assign _T_92742 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[LoadQueue.scala 238:96:@38272.8]
  assign _T_92750 = {lastConflict_5_15,lastConflict_5_14,lastConflict_5_13,lastConflict_5_12,lastConflict_5_11,lastConflict_5_10,lastConflict_5_9,lastConflict_5_8,_T_92742}; // @[LoadQueue.scala 238:96:@38280.8]
  assign _T_92751 = _T_92735 < _T_92750; // @[LoadQueue.scala 238:61:@38281.8]
  assign _T_92752 = canBypass_5 & _T_92751; // @[LoadQueue.scala 237:64:@38282.8]
  assign _GEN_1989 = _T_92681 ? _T_92752 : 1'h0; // @[LoadQueue.scala 230:110:@38214.6]
  assign bypassRequest_5 = _T_92673 ? _GEN_1989 : 1'h0; // @[LoadQueue.scala 229:71:@38208.4]
  assign _GEN_1946 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[LoadQueue.scala 217:34:@37721.6]
  assign _GEN_1947 = initBits_5 ? 1'h0 : _GEN_1946; // @[LoadQueue.scala 215:23:@37717.4]
  assign _T_92811 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[LoadQueue.scala 238:58:@38339.8]
  assign _T_92819 = {storeAddrNotKnownFlagsPReg_6_15,storeAddrNotKnownFlagsPReg_6_14,storeAddrNotKnownFlagsPReg_6_13,storeAddrNotKnownFlagsPReg_6_12,storeAddrNotKnownFlagsPReg_6_11,storeAddrNotKnownFlagsPReg_6_10,storeAddrNotKnownFlagsPReg_6_9,storeAddrNotKnownFlagsPReg_6_8,_T_92811}; // @[LoadQueue.scala 238:58:@38347.8]
  assign _T_92826 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[LoadQueue.scala 238:96:@38354.8]
  assign _T_92834 = {lastConflict_6_15,lastConflict_6_14,lastConflict_6_13,lastConflict_6_12,lastConflict_6_11,lastConflict_6_10,lastConflict_6_9,lastConflict_6_8,_T_92826}; // @[LoadQueue.scala 238:96:@38362.8]
  assign _T_92835 = _T_92819 < _T_92834; // @[LoadQueue.scala 238:61:@38363.8]
  assign _T_92836 = canBypass_6 & _T_92835; // @[LoadQueue.scala 237:64:@38364.8]
  assign _GEN_1993 = _T_92765 ? _T_92836 : 1'h0; // @[LoadQueue.scala 230:110:@38296.6]
  assign bypassRequest_6 = _T_92757 ? _GEN_1993 : 1'h0; // @[LoadQueue.scala 229:71:@38290.4]
  assign _GEN_1948 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[LoadQueue.scala 217:34:@37728.6]
  assign _GEN_1949 = initBits_6 ? 1'h0 : _GEN_1948; // @[LoadQueue.scala 215:23:@37724.4]
  assign _T_92895 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[LoadQueue.scala 238:58:@38421.8]
  assign _T_92903 = {storeAddrNotKnownFlagsPReg_7_15,storeAddrNotKnownFlagsPReg_7_14,storeAddrNotKnownFlagsPReg_7_13,storeAddrNotKnownFlagsPReg_7_12,storeAddrNotKnownFlagsPReg_7_11,storeAddrNotKnownFlagsPReg_7_10,storeAddrNotKnownFlagsPReg_7_9,storeAddrNotKnownFlagsPReg_7_8,_T_92895}; // @[LoadQueue.scala 238:58:@38429.8]
  assign _T_92910 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[LoadQueue.scala 238:96:@38436.8]
  assign _T_92918 = {lastConflict_7_15,lastConflict_7_14,lastConflict_7_13,lastConflict_7_12,lastConflict_7_11,lastConflict_7_10,lastConflict_7_9,lastConflict_7_8,_T_92910}; // @[LoadQueue.scala 238:96:@38444.8]
  assign _T_92919 = _T_92903 < _T_92918; // @[LoadQueue.scala 238:61:@38445.8]
  assign _T_92920 = canBypass_7 & _T_92919; // @[LoadQueue.scala 237:64:@38446.8]
  assign _GEN_1997 = _T_92849 ? _T_92920 : 1'h0; // @[LoadQueue.scala 230:110:@38378.6]
  assign bypassRequest_7 = _T_92841 ? _GEN_1997 : 1'h0; // @[LoadQueue.scala 229:71:@38372.4]
  assign _GEN_1950 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[LoadQueue.scala 217:34:@37735.6]
  assign _GEN_1951 = initBits_7 ? 1'h0 : _GEN_1950; // @[LoadQueue.scala 215:23:@37731.4]
  assign _T_92979 = {storeAddrNotKnownFlagsPReg_8_7,storeAddrNotKnownFlagsPReg_8_6,storeAddrNotKnownFlagsPReg_8_5,storeAddrNotKnownFlagsPReg_8_4,storeAddrNotKnownFlagsPReg_8_3,storeAddrNotKnownFlagsPReg_8_2,storeAddrNotKnownFlagsPReg_8_1,storeAddrNotKnownFlagsPReg_8_0}; // @[LoadQueue.scala 238:58:@38503.8]
  assign _T_92987 = {storeAddrNotKnownFlagsPReg_8_15,storeAddrNotKnownFlagsPReg_8_14,storeAddrNotKnownFlagsPReg_8_13,storeAddrNotKnownFlagsPReg_8_12,storeAddrNotKnownFlagsPReg_8_11,storeAddrNotKnownFlagsPReg_8_10,storeAddrNotKnownFlagsPReg_8_9,storeAddrNotKnownFlagsPReg_8_8,_T_92979}; // @[LoadQueue.scala 238:58:@38511.8]
  assign _T_92994 = {lastConflict_8_7,lastConflict_8_6,lastConflict_8_5,lastConflict_8_4,lastConflict_8_3,lastConflict_8_2,lastConflict_8_1,lastConflict_8_0}; // @[LoadQueue.scala 238:96:@38518.8]
  assign _T_93002 = {lastConflict_8_15,lastConflict_8_14,lastConflict_8_13,lastConflict_8_12,lastConflict_8_11,lastConflict_8_10,lastConflict_8_9,lastConflict_8_8,_T_92994}; // @[LoadQueue.scala 238:96:@38526.8]
  assign _T_93003 = _T_92987 < _T_93002; // @[LoadQueue.scala 238:61:@38527.8]
  assign _T_93004 = canBypass_8 & _T_93003; // @[LoadQueue.scala 237:64:@38528.8]
  assign _GEN_2001 = _T_92933 ? _T_93004 : 1'h0; // @[LoadQueue.scala 230:110:@38460.6]
  assign bypassRequest_8 = _T_92925 ? _GEN_2001 : 1'h0; // @[LoadQueue.scala 229:71:@38454.4]
  assign _GEN_1952 = bypassRequest_8 ? 1'h1 : bypassInitiated_8; // @[LoadQueue.scala 217:34:@37742.6]
  assign _GEN_1953 = initBits_8 ? 1'h0 : _GEN_1952; // @[LoadQueue.scala 215:23:@37738.4]
  assign _T_93063 = {storeAddrNotKnownFlagsPReg_9_7,storeAddrNotKnownFlagsPReg_9_6,storeAddrNotKnownFlagsPReg_9_5,storeAddrNotKnownFlagsPReg_9_4,storeAddrNotKnownFlagsPReg_9_3,storeAddrNotKnownFlagsPReg_9_2,storeAddrNotKnownFlagsPReg_9_1,storeAddrNotKnownFlagsPReg_9_0}; // @[LoadQueue.scala 238:58:@38585.8]
  assign _T_93071 = {storeAddrNotKnownFlagsPReg_9_15,storeAddrNotKnownFlagsPReg_9_14,storeAddrNotKnownFlagsPReg_9_13,storeAddrNotKnownFlagsPReg_9_12,storeAddrNotKnownFlagsPReg_9_11,storeAddrNotKnownFlagsPReg_9_10,storeAddrNotKnownFlagsPReg_9_9,storeAddrNotKnownFlagsPReg_9_8,_T_93063}; // @[LoadQueue.scala 238:58:@38593.8]
  assign _T_93078 = {lastConflict_9_7,lastConflict_9_6,lastConflict_9_5,lastConflict_9_4,lastConflict_9_3,lastConflict_9_2,lastConflict_9_1,lastConflict_9_0}; // @[LoadQueue.scala 238:96:@38600.8]
  assign _T_93086 = {lastConflict_9_15,lastConflict_9_14,lastConflict_9_13,lastConflict_9_12,lastConflict_9_11,lastConflict_9_10,lastConflict_9_9,lastConflict_9_8,_T_93078}; // @[LoadQueue.scala 238:96:@38608.8]
  assign _T_93087 = _T_93071 < _T_93086; // @[LoadQueue.scala 238:61:@38609.8]
  assign _T_93088 = canBypass_9 & _T_93087; // @[LoadQueue.scala 237:64:@38610.8]
  assign _GEN_2005 = _T_93017 ? _T_93088 : 1'h0; // @[LoadQueue.scala 230:110:@38542.6]
  assign bypassRequest_9 = _T_93009 ? _GEN_2005 : 1'h0; // @[LoadQueue.scala 229:71:@38536.4]
  assign _GEN_1954 = bypassRequest_9 ? 1'h1 : bypassInitiated_9; // @[LoadQueue.scala 217:34:@37749.6]
  assign _GEN_1955 = initBits_9 ? 1'h0 : _GEN_1954; // @[LoadQueue.scala 215:23:@37745.4]
  assign _T_93147 = {storeAddrNotKnownFlagsPReg_10_7,storeAddrNotKnownFlagsPReg_10_6,storeAddrNotKnownFlagsPReg_10_5,storeAddrNotKnownFlagsPReg_10_4,storeAddrNotKnownFlagsPReg_10_3,storeAddrNotKnownFlagsPReg_10_2,storeAddrNotKnownFlagsPReg_10_1,storeAddrNotKnownFlagsPReg_10_0}; // @[LoadQueue.scala 238:58:@38667.8]
  assign _T_93155 = {storeAddrNotKnownFlagsPReg_10_15,storeAddrNotKnownFlagsPReg_10_14,storeAddrNotKnownFlagsPReg_10_13,storeAddrNotKnownFlagsPReg_10_12,storeAddrNotKnownFlagsPReg_10_11,storeAddrNotKnownFlagsPReg_10_10,storeAddrNotKnownFlagsPReg_10_9,storeAddrNotKnownFlagsPReg_10_8,_T_93147}; // @[LoadQueue.scala 238:58:@38675.8]
  assign _T_93162 = {lastConflict_10_7,lastConflict_10_6,lastConflict_10_5,lastConflict_10_4,lastConflict_10_3,lastConflict_10_2,lastConflict_10_1,lastConflict_10_0}; // @[LoadQueue.scala 238:96:@38682.8]
  assign _T_93170 = {lastConflict_10_15,lastConflict_10_14,lastConflict_10_13,lastConflict_10_12,lastConflict_10_11,lastConflict_10_10,lastConflict_10_9,lastConflict_10_8,_T_93162}; // @[LoadQueue.scala 238:96:@38690.8]
  assign _T_93171 = _T_93155 < _T_93170; // @[LoadQueue.scala 238:61:@38691.8]
  assign _T_93172 = canBypass_10 & _T_93171; // @[LoadQueue.scala 237:64:@38692.8]
  assign _GEN_2009 = _T_93101 ? _T_93172 : 1'h0; // @[LoadQueue.scala 230:110:@38624.6]
  assign bypassRequest_10 = _T_93093 ? _GEN_2009 : 1'h0; // @[LoadQueue.scala 229:71:@38618.4]
  assign _GEN_1956 = bypassRequest_10 ? 1'h1 : bypassInitiated_10; // @[LoadQueue.scala 217:34:@37756.6]
  assign _GEN_1957 = initBits_10 ? 1'h0 : _GEN_1956; // @[LoadQueue.scala 215:23:@37752.4]
  assign _T_93231 = {storeAddrNotKnownFlagsPReg_11_7,storeAddrNotKnownFlagsPReg_11_6,storeAddrNotKnownFlagsPReg_11_5,storeAddrNotKnownFlagsPReg_11_4,storeAddrNotKnownFlagsPReg_11_3,storeAddrNotKnownFlagsPReg_11_2,storeAddrNotKnownFlagsPReg_11_1,storeAddrNotKnownFlagsPReg_11_0}; // @[LoadQueue.scala 238:58:@38749.8]
  assign _T_93239 = {storeAddrNotKnownFlagsPReg_11_15,storeAddrNotKnownFlagsPReg_11_14,storeAddrNotKnownFlagsPReg_11_13,storeAddrNotKnownFlagsPReg_11_12,storeAddrNotKnownFlagsPReg_11_11,storeAddrNotKnownFlagsPReg_11_10,storeAddrNotKnownFlagsPReg_11_9,storeAddrNotKnownFlagsPReg_11_8,_T_93231}; // @[LoadQueue.scala 238:58:@38757.8]
  assign _T_93246 = {lastConflict_11_7,lastConflict_11_6,lastConflict_11_5,lastConflict_11_4,lastConflict_11_3,lastConflict_11_2,lastConflict_11_1,lastConflict_11_0}; // @[LoadQueue.scala 238:96:@38764.8]
  assign _T_93254 = {lastConflict_11_15,lastConflict_11_14,lastConflict_11_13,lastConflict_11_12,lastConflict_11_11,lastConflict_11_10,lastConflict_11_9,lastConflict_11_8,_T_93246}; // @[LoadQueue.scala 238:96:@38772.8]
  assign _T_93255 = _T_93239 < _T_93254; // @[LoadQueue.scala 238:61:@38773.8]
  assign _T_93256 = canBypass_11 & _T_93255; // @[LoadQueue.scala 237:64:@38774.8]
  assign _GEN_2013 = _T_93185 ? _T_93256 : 1'h0; // @[LoadQueue.scala 230:110:@38706.6]
  assign bypassRequest_11 = _T_93177 ? _GEN_2013 : 1'h0; // @[LoadQueue.scala 229:71:@38700.4]
  assign _GEN_1958 = bypassRequest_11 ? 1'h1 : bypassInitiated_11; // @[LoadQueue.scala 217:34:@37763.6]
  assign _GEN_1959 = initBits_11 ? 1'h0 : _GEN_1958; // @[LoadQueue.scala 215:23:@37759.4]
  assign _T_93315 = {storeAddrNotKnownFlagsPReg_12_7,storeAddrNotKnownFlagsPReg_12_6,storeAddrNotKnownFlagsPReg_12_5,storeAddrNotKnownFlagsPReg_12_4,storeAddrNotKnownFlagsPReg_12_3,storeAddrNotKnownFlagsPReg_12_2,storeAddrNotKnownFlagsPReg_12_1,storeAddrNotKnownFlagsPReg_12_0}; // @[LoadQueue.scala 238:58:@38831.8]
  assign _T_93323 = {storeAddrNotKnownFlagsPReg_12_15,storeAddrNotKnownFlagsPReg_12_14,storeAddrNotKnownFlagsPReg_12_13,storeAddrNotKnownFlagsPReg_12_12,storeAddrNotKnownFlagsPReg_12_11,storeAddrNotKnownFlagsPReg_12_10,storeAddrNotKnownFlagsPReg_12_9,storeAddrNotKnownFlagsPReg_12_8,_T_93315}; // @[LoadQueue.scala 238:58:@38839.8]
  assign _T_93330 = {lastConflict_12_7,lastConflict_12_6,lastConflict_12_5,lastConflict_12_4,lastConflict_12_3,lastConflict_12_2,lastConflict_12_1,lastConflict_12_0}; // @[LoadQueue.scala 238:96:@38846.8]
  assign _T_93338 = {lastConflict_12_15,lastConflict_12_14,lastConflict_12_13,lastConflict_12_12,lastConflict_12_11,lastConflict_12_10,lastConflict_12_9,lastConflict_12_8,_T_93330}; // @[LoadQueue.scala 238:96:@38854.8]
  assign _T_93339 = _T_93323 < _T_93338; // @[LoadQueue.scala 238:61:@38855.8]
  assign _T_93340 = canBypass_12 & _T_93339; // @[LoadQueue.scala 237:64:@38856.8]
  assign _GEN_2017 = _T_93269 ? _T_93340 : 1'h0; // @[LoadQueue.scala 230:110:@38788.6]
  assign bypassRequest_12 = _T_93261 ? _GEN_2017 : 1'h0; // @[LoadQueue.scala 229:71:@38782.4]
  assign _GEN_1960 = bypassRequest_12 ? 1'h1 : bypassInitiated_12; // @[LoadQueue.scala 217:34:@37770.6]
  assign _GEN_1961 = initBits_12 ? 1'h0 : _GEN_1960; // @[LoadQueue.scala 215:23:@37766.4]
  assign _T_93399 = {storeAddrNotKnownFlagsPReg_13_7,storeAddrNotKnownFlagsPReg_13_6,storeAddrNotKnownFlagsPReg_13_5,storeAddrNotKnownFlagsPReg_13_4,storeAddrNotKnownFlagsPReg_13_3,storeAddrNotKnownFlagsPReg_13_2,storeAddrNotKnownFlagsPReg_13_1,storeAddrNotKnownFlagsPReg_13_0}; // @[LoadQueue.scala 238:58:@38913.8]
  assign _T_93407 = {storeAddrNotKnownFlagsPReg_13_15,storeAddrNotKnownFlagsPReg_13_14,storeAddrNotKnownFlagsPReg_13_13,storeAddrNotKnownFlagsPReg_13_12,storeAddrNotKnownFlagsPReg_13_11,storeAddrNotKnownFlagsPReg_13_10,storeAddrNotKnownFlagsPReg_13_9,storeAddrNotKnownFlagsPReg_13_8,_T_93399}; // @[LoadQueue.scala 238:58:@38921.8]
  assign _T_93414 = {lastConflict_13_7,lastConflict_13_6,lastConflict_13_5,lastConflict_13_4,lastConflict_13_3,lastConflict_13_2,lastConflict_13_1,lastConflict_13_0}; // @[LoadQueue.scala 238:96:@38928.8]
  assign _T_93422 = {lastConflict_13_15,lastConflict_13_14,lastConflict_13_13,lastConflict_13_12,lastConflict_13_11,lastConflict_13_10,lastConflict_13_9,lastConflict_13_8,_T_93414}; // @[LoadQueue.scala 238:96:@38936.8]
  assign _T_93423 = _T_93407 < _T_93422; // @[LoadQueue.scala 238:61:@38937.8]
  assign _T_93424 = canBypass_13 & _T_93423; // @[LoadQueue.scala 237:64:@38938.8]
  assign _GEN_2021 = _T_93353 ? _T_93424 : 1'h0; // @[LoadQueue.scala 230:110:@38870.6]
  assign bypassRequest_13 = _T_93345 ? _GEN_2021 : 1'h0; // @[LoadQueue.scala 229:71:@38864.4]
  assign _GEN_1962 = bypassRequest_13 ? 1'h1 : bypassInitiated_13; // @[LoadQueue.scala 217:34:@37777.6]
  assign _GEN_1963 = initBits_13 ? 1'h0 : _GEN_1962; // @[LoadQueue.scala 215:23:@37773.4]
  assign _T_93483 = {storeAddrNotKnownFlagsPReg_14_7,storeAddrNotKnownFlagsPReg_14_6,storeAddrNotKnownFlagsPReg_14_5,storeAddrNotKnownFlagsPReg_14_4,storeAddrNotKnownFlagsPReg_14_3,storeAddrNotKnownFlagsPReg_14_2,storeAddrNotKnownFlagsPReg_14_1,storeAddrNotKnownFlagsPReg_14_0}; // @[LoadQueue.scala 238:58:@38995.8]
  assign _T_93491 = {storeAddrNotKnownFlagsPReg_14_15,storeAddrNotKnownFlagsPReg_14_14,storeAddrNotKnownFlagsPReg_14_13,storeAddrNotKnownFlagsPReg_14_12,storeAddrNotKnownFlagsPReg_14_11,storeAddrNotKnownFlagsPReg_14_10,storeAddrNotKnownFlagsPReg_14_9,storeAddrNotKnownFlagsPReg_14_8,_T_93483}; // @[LoadQueue.scala 238:58:@39003.8]
  assign _T_93498 = {lastConflict_14_7,lastConflict_14_6,lastConflict_14_5,lastConflict_14_4,lastConflict_14_3,lastConflict_14_2,lastConflict_14_1,lastConflict_14_0}; // @[LoadQueue.scala 238:96:@39010.8]
  assign _T_93506 = {lastConflict_14_15,lastConflict_14_14,lastConflict_14_13,lastConflict_14_12,lastConflict_14_11,lastConflict_14_10,lastConflict_14_9,lastConflict_14_8,_T_93498}; // @[LoadQueue.scala 238:96:@39018.8]
  assign _T_93507 = _T_93491 < _T_93506; // @[LoadQueue.scala 238:61:@39019.8]
  assign _T_93508 = canBypass_14 & _T_93507; // @[LoadQueue.scala 237:64:@39020.8]
  assign _GEN_2025 = _T_93437 ? _T_93508 : 1'h0; // @[LoadQueue.scala 230:110:@38952.6]
  assign bypassRequest_14 = _T_93429 ? _GEN_2025 : 1'h0; // @[LoadQueue.scala 229:71:@38946.4]
  assign _GEN_1964 = bypassRequest_14 ? 1'h1 : bypassInitiated_14; // @[LoadQueue.scala 217:34:@37784.6]
  assign _GEN_1965 = initBits_14 ? 1'h0 : _GEN_1964; // @[LoadQueue.scala 215:23:@37780.4]
  assign _T_93567 = {storeAddrNotKnownFlagsPReg_15_7,storeAddrNotKnownFlagsPReg_15_6,storeAddrNotKnownFlagsPReg_15_5,storeAddrNotKnownFlagsPReg_15_4,storeAddrNotKnownFlagsPReg_15_3,storeAddrNotKnownFlagsPReg_15_2,storeAddrNotKnownFlagsPReg_15_1,storeAddrNotKnownFlagsPReg_15_0}; // @[LoadQueue.scala 238:58:@39077.8]
  assign _T_93575 = {storeAddrNotKnownFlagsPReg_15_15,storeAddrNotKnownFlagsPReg_15_14,storeAddrNotKnownFlagsPReg_15_13,storeAddrNotKnownFlagsPReg_15_12,storeAddrNotKnownFlagsPReg_15_11,storeAddrNotKnownFlagsPReg_15_10,storeAddrNotKnownFlagsPReg_15_9,storeAddrNotKnownFlagsPReg_15_8,_T_93567}; // @[LoadQueue.scala 238:58:@39085.8]
  assign _T_93582 = {lastConflict_15_7,lastConflict_15_6,lastConflict_15_5,lastConflict_15_4,lastConflict_15_3,lastConflict_15_2,lastConflict_15_1,lastConflict_15_0}; // @[LoadQueue.scala 238:96:@39092.8]
  assign _T_93590 = {lastConflict_15_15,lastConflict_15_14,lastConflict_15_13,lastConflict_15_12,lastConflict_15_11,lastConflict_15_10,lastConflict_15_9,lastConflict_15_8,_T_93582}; // @[LoadQueue.scala 238:96:@39100.8]
  assign _T_93591 = _T_93575 < _T_93590; // @[LoadQueue.scala 238:61:@39101.8]
  assign _T_93592 = canBypass_15 & _T_93591; // @[LoadQueue.scala 237:64:@39102.8]
  assign _GEN_2029 = _T_93521 ? _T_93592 : 1'h0; // @[LoadQueue.scala 230:110:@39034.6]
  assign bypassRequest_15 = _T_93513 ? _GEN_2029 : 1'h0; // @[LoadQueue.scala 229:71:@39028.4]
  assign _GEN_1966 = bypassRequest_15 ? 1'h1 : bypassInitiated_15; // @[LoadQueue.scala 217:34:@37791.6]
  assign _GEN_1967 = initBits_15 ? 1'h0 : _GEN_1966; // @[LoadQueue.scala 215:23:@37787.4]
  assign _T_93596 = loadRequest_0 | loadRequest_1; // @[LoadQueue.scala 247:28:@39108.4]
  assign _T_93597 = _T_93596 | loadRequest_2; // @[LoadQueue.scala 247:28:@39109.4]
  assign _T_93598 = _T_93597 | loadRequest_3; // @[LoadQueue.scala 247:28:@39110.4]
  assign _T_93599 = _T_93598 | loadRequest_4; // @[LoadQueue.scala 247:28:@39111.4]
  assign _T_93600 = _T_93599 | loadRequest_5; // @[LoadQueue.scala 247:28:@39112.4]
  assign _T_93601 = _T_93600 | loadRequest_6; // @[LoadQueue.scala 247:28:@39113.4]
  assign _T_93602 = _T_93601 | loadRequest_7; // @[LoadQueue.scala 247:28:@39114.4]
  assign _T_93603 = _T_93602 | loadRequest_8; // @[LoadQueue.scala 247:28:@39115.4]
  assign _T_93604 = _T_93603 | loadRequest_9; // @[LoadQueue.scala 247:28:@39116.4]
  assign _T_93605 = _T_93604 | loadRequest_10; // @[LoadQueue.scala 247:28:@39117.4]
  assign _T_93606 = _T_93605 | loadRequest_11; // @[LoadQueue.scala 247:28:@39118.4]
  assign _T_93607 = _T_93606 | loadRequest_12; // @[LoadQueue.scala 247:28:@39119.4]
  assign _T_93608 = _T_93607 | loadRequest_13; // @[LoadQueue.scala 247:28:@39120.4]
  assign _T_93609 = _T_93608 | loadRequest_14; // @[LoadQueue.scala 247:28:@39121.4]
  assign _T_93610 = _T_93609 | loadRequest_15; // @[LoadQueue.scala 247:28:@39122.4]
  assign _T_93627 = priorityLoadRequest_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@39124.6]
  assign _T_93628 = priorityLoadRequest_13 ? 4'hd : _T_93627; // @[Mux.scala 31:69:@39125.6]
  assign _T_93629 = priorityLoadRequest_12 ? 4'hc : _T_93628; // @[Mux.scala 31:69:@39126.6]
  assign _T_93630 = priorityLoadRequest_11 ? 4'hb : _T_93629; // @[Mux.scala 31:69:@39127.6]
  assign _T_93631 = priorityLoadRequest_10 ? 4'ha : _T_93630; // @[Mux.scala 31:69:@39128.6]
  assign _T_93632 = priorityLoadRequest_9 ? 4'h9 : _T_93631; // @[Mux.scala 31:69:@39129.6]
  assign _T_93633 = priorityLoadRequest_8 ? 4'h8 : _T_93632; // @[Mux.scala 31:69:@39130.6]
  assign _T_93634 = priorityLoadRequest_7 ? 4'h7 : _T_93633; // @[Mux.scala 31:69:@39131.6]
  assign _T_93635 = priorityLoadRequest_6 ? 4'h6 : _T_93634; // @[Mux.scala 31:69:@39132.6]
  assign _T_93636 = priorityLoadRequest_5 ? 4'h5 : _T_93635; // @[Mux.scala 31:69:@39133.6]
  assign _T_93637 = priorityLoadRequest_4 ? 4'h4 : _T_93636; // @[Mux.scala 31:69:@39134.6]
  assign _T_93638 = priorityLoadRequest_3 ? 4'h3 : _T_93637; // @[Mux.scala 31:69:@39135.6]
  assign _T_93639 = priorityLoadRequest_2 ? 4'h2 : _T_93638; // @[Mux.scala 31:69:@39136.6]
  assign _T_93640 = priorityLoadRequest_1 ? 4'h1 : _T_93639; // @[Mux.scala 31:69:@39137.6]
  assign _T_93641 = priorityLoadRequest_0 ? 4'h0 : _T_93640; // @[Mux.scala 31:69:@39138.6]
  assign _GEN_2033 = 4'h1 == _T_93641 ? addrQ_1 : addrQ_0; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2034 = 4'h2 == _T_93641 ? addrQ_2 : _GEN_2033; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2035 = 4'h3 == _T_93641 ? addrQ_3 : _GEN_2034; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2036 = 4'h4 == _T_93641 ? addrQ_4 : _GEN_2035; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2037 = 4'h5 == _T_93641 ? addrQ_5 : _GEN_2036; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2038 = 4'h6 == _T_93641 ? addrQ_6 : _GEN_2037; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2039 = 4'h7 == _T_93641 ? addrQ_7 : _GEN_2038; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2040 = 4'h8 == _T_93641 ? addrQ_8 : _GEN_2039; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2041 = 4'h9 == _T_93641 ? addrQ_9 : _GEN_2040; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2042 = 4'ha == _T_93641 ? addrQ_10 : _GEN_2041; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2043 = 4'hb == _T_93641 ? addrQ_11 : _GEN_2042; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2044 = 4'hc == _T_93641 ? addrQ_12 : _GEN_2043; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2045 = 4'hd == _T_93641 ? addrQ_13 : _GEN_2044; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2046 = 4'he == _T_93641 ? addrQ_14 : _GEN_2045; // @[LoadQueue.scala 248:24:@39139.6]
  assign _GEN_2047 = 4'hf == _T_93641 ? addrQ_15 : _GEN_2046; // @[LoadQueue.scala 248:24:@39139.6]
  assign _T_93649 = prevPriorityRequest_0 | bypassRequest_0; // @[LoadQueue.scala 261:41:@39150.6]
  assign _GEN_2050 = _T_93649 ? 1'h1 : dataKnown_0; // @[LoadQueue.scala 261:62:@39151.6]
  assign _GEN_2051 = initBits_0 ? 1'h0 : _GEN_2050; // @[LoadQueue.scala 259:25:@39146.4]
  assign _T_93652 = prevPriorityRequest_1 | bypassRequest_1; // @[LoadQueue.scala 261:41:@39158.6]
  assign _GEN_2052 = _T_93652 ? 1'h1 : dataKnown_1; // @[LoadQueue.scala 261:62:@39159.6]
  assign _GEN_2053 = initBits_1 ? 1'h0 : _GEN_2052; // @[LoadQueue.scala 259:25:@39154.4]
  assign _T_93655 = prevPriorityRequest_2 | bypassRequest_2; // @[LoadQueue.scala 261:41:@39166.6]
  assign _GEN_2054 = _T_93655 ? 1'h1 : dataKnown_2; // @[LoadQueue.scala 261:62:@39167.6]
  assign _GEN_2055 = initBits_2 ? 1'h0 : _GEN_2054; // @[LoadQueue.scala 259:25:@39162.4]
  assign _T_93658 = prevPriorityRequest_3 | bypassRequest_3; // @[LoadQueue.scala 261:41:@39174.6]
  assign _GEN_2056 = _T_93658 ? 1'h1 : dataKnown_3; // @[LoadQueue.scala 261:62:@39175.6]
  assign _GEN_2057 = initBits_3 ? 1'h0 : _GEN_2056; // @[LoadQueue.scala 259:25:@39170.4]
  assign _T_93661 = prevPriorityRequest_4 | bypassRequest_4; // @[LoadQueue.scala 261:41:@39182.6]
  assign _GEN_2058 = _T_93661 ? 1'h1 : dataKnown_4; // @[LoadQueue.scala 261:62:@39183.6]
  assign _GEN_2059 = initBits_4 ? 1'h0 : _GEN_2058; // @[LoadQueue.scala 259:25:@39178.4]
  assign _T_93664 = prevPriorityRequest_5 | bypassRequest_5; // @[LoadQueue.scala 261:41:@39190.6]
  assign _GEN_2060 = _T_93664 ? 1'h1 : dataKnown_5; // @[LoadQueue.scala 261:62:@39191.6]
  assign _GEN_2061 = initBits_5 ? 1'h0 : _GEN_2060; // @[LoadQueue.scala 259:25:@39186.4]
  assign _T_93667 = prevPriorityRequest_6 | bypassRequest_6; // @[LoadQueue.scala 261:41:@39198.6]
  assign _GEN_2062 = _T_93667 ? 1'h1 : dataKnown_6; // @[LoadQueue.scala 261:62:@39199.6]
  assign _GEN_2063 = initBits_6 ? 1'h0 : _GEN_2062; // @[LoadQueue.scala 259:25:@39194.4]
  assign _T_93670 = prevPriorityRequest_7 | bypassRequest_7; // @[LoadQueue.scala 261:41:@39206.6]
  assign _GEN_2064 = _T_93670 ? 1'h1 : dataKnown_7; // @[LoadQueue.scala 261:62:@39207.6]
  assign _GEN_2065 = initBits_7 ? 1'h0 : _GEN_2064; // @[LoadQueue.scala 259:25:@39202.4]
  assign _T_93673 = prevPriorityRequest_8 | bypassRequest_8; // @[LoadQueue.scala 261:41:@39214.6]
  assign _GEN_2066 = _T_93673 ? 1'h1 : dataKnown_8; // @[LoadQueue.scala 261:62:@39215.6]
  assign _GEN_2067 = initBits_8 ? 1'h0 : _GEN_2066; // @[LoadQueue.scala 259:25:@39210.4]
  assign _T_93676 = prevPriorityRequest_9 | bypassRequest_9; // @[LoadQueue.scala 261:41:@39222.6]
  assign _GEN_2068 = _T_93676 ? 1'h1 : dataKnown_9; // @[LoadQueue.scala 261:62:@39223.6]
  assign _GEN_2069 = initBits_9 ? 1'h0 : _GEN_2068; // @[LoadQueue.scala 259:25:@39218.4]
  assign _T_93679 = prevPriorityRequest_10 | bypassRequest_10; // @[LoadQueue.scala 261:41:@39230.6]
  assign _GEN_2070 = _T_93679 ? 1'h1 : dataKnown_10; // @[LoadQueue.scala 261:62:@39231.6]
  assign _GEN_2071 = initBits_10 ? 1'h0 : _GEN_2070; // @[LoadQueue.scala 259:25:@39226.4]
  assign _T_93682 = prevPriorityRequest_11 | bypassRequest_11; // @[LoadQueue.scala 261:41:@39238.6]
  assign _GEN_2072 = _T_93682 ? 1'h1 : dataKnown_11; // @[LoadQueue.scala 261:62:@39239.6]
  assign _GEN_2073 = initBits_11 ? 1'h0 : _GEN_2072; // @[LoadQueue.scala 259:25:@39234.4]
  assign _T_93685 = prevPriorityRequest_12 | bypassRequest_12; // @[LoadQueue.scala 261:41:@39246.6]
  assign _GEN_2074 = _T_93685 ? 1'h1 : dataKnown_12; // @[LoadQueue.scala 261:62:@39247.6]
  assign _GEN_2075 = initBits_12 ? 1'h0 : _GEN_2074; // @[LoadQueue.scala 259:25:@39242.4]
  assign _T_93688 = prevPriorityRequest_13 | bypassRequest_13; // @[LoadQueue.scala 261:41:@39254.6]
  assign _GEN_2076 = _T_93688 ? 1'h1 : dataKnown_13; // @[LoadQueue.scala 261:62:@39255.6]
  assign _GEN_2077 = initBits_13 ? 1'h0 : _GEN_2076; // @[LoadQueue.scala 259:25:@39250.4]
  assign _T_93691 = prevPriorityRequest_14 | bypassRequest_14; // @[LoadQueue.scala 261:41:@39262.6]
  assign _GEN_2078 = _T_93691 ? 1'h1 : dataKnown_14; // @[LoadQueue.scala 261:62:@39263.6]
  assign _GEN_2079 = initBits_14 ? 1'h0 : _GEN_2078; // @[LoadQueue.scala 259:25:@39258.4]
  assign _T_93694 = prevPriorityRequest_15 | bypassRequest_15; // @[LoadQueue.scala 261:41:@39270.6]
  assign _GEN_2080 = _T_93694 ? 1'h1 : dataKnown_15; // @[LoadQueue.scala 261:62:@39271.6]
  assign _GEN_2081 = initBits_15 ? 1'h0 : _GEN_2080; // @[LoadQueue.scala 259:25:@39266.4]
  assign _GEN_2082 = prevPriorityRequest_0 ? io_loadDataFromMem : dataQ_0; // @[LoadQueue.scala 269:44:@39278.6]
  assign _GEN_2083 = bypassRequest_0 ? bypassVal_0 : _GEN_2082; // @[LoadQueue.scala 267:32:@39274.4]
  assign _GEN_2084 = prevPriorityRequest_1 ? io_loadDataFromMem : dataQ_1; // @[LoadQueue.scala 269:44:@39285.6]
  assign _GEN_2085 = bypassRequest_1 ? bypassVal_1 : _GEN_2084; // @[LoadQueue.scala 267:32:@39281.4]
  assign _GEN_2086 = prevPriorityRequest_2 ? io_loadDataFromMem : dataQ_2; // @[LoadQueue.scala 269:44:@39292.6]
  assign _GEN_2087 = bypassRequest_2 ? bypassVal_2 : _GEN_2086; // @[LoadQueue.scala 267:32:@39288.4]
  assign _GEN_2088 = prevPriorityRequest_3 ? io_loadDataFromMem : dataQ_3; // @[LoadQueue.scala 269:44:@39299.6]
  assign _GEN_2089 = bypassRequest_3 ? bypassVal_3 : _GEN_2088; // @[LoadQueue.scala 267:32:@39295.4]
  assign _GEN_2090 = prevPriorityRequest_4 ? io_loadDataFromMem : dataQ_4; // @[LoadQueue.scala 269:44:@39306.6]
  assign _GEN_2091 = bypassRequest_4 ? bypassVal_4 : _GEN_2090; // @[LoadQueue.scala 267:32:@39302.4]
  assign _GEN_2092 = prevPriorityRequest_5 ? io_loadDataFromMem : dataQ_5; // @[LoadQueue.scala 269:44:@39313.6]
  assign _GEN_2093 = bypassRequest_5 ? bypassVal_5 : _GEN_2092; // @[LoadQueue.scala 267:32:@39309.4]
  assign _GEN_2094 = prevPriorityRequest_6 ? io_loadDataFromMem : dataQ_6; // @[LoadQueue.scala 269:44:@39320.6]
  assign _GEN_2095 = bypassRequest_6 ? bypassVal_6 : _GEN_2094; // @[LoadQueue.scala 267:32:@39316.4]
  assign _GEN_2096 = prevPriorityRequest_7 ? io_loadDataFromMem : dataQ_7; // @[LoadQueue.scala 269:44:@39327.6]
  assign _GEN_2097 = bypassRequest_7 ? bypassVal_7 : _GEN_2096; // @[LoadQueue.scala 267:32:@39323.4]
  assign _GEN_2098 = prevPriorityRequest_8 ? io_loadDataFromMem : dataQ_8; // @[LoadQueue.scala 269:44:@39334.6]
  assign _GEN_2099 = bypassRequest_8 ? bypassVal_8 : _GEN_2098; // @[LoadQueue.scala 267:32:@39330.4]
  assign _GEN_2100 = prevPriorityRequest_9 ? io_loadDataFromMem : dataQ_9; // @[LoadQueue.scala 269:44:@39341.6]
  assign _GEN_2101 = bypassRequest_9 ? bypassVal_9 : _GEN_2100; // @[LoadQueue.scala 267:32:@39337.4]
  assign _GEN_2102 = prevPriorityRequest_10 ? io_loadDataFromMem : dataQ_10; // @[LoadQueue.scala 269:44:@39348.6]
  assign _GEN_2103 = bypassRequest_10 ? bypassVal_10 : _GEN_2102; // @[LoadQueue.scala 267:32:@39344.4]
  assign _GEN_2104 = prevPriorityRequest_11 ? io_loadDataFromMem : dataQ_11; // @[LoadQueue.scala 269:44:@39355.6]
  assign _GEN_2105 = bypassRequest_11 ? bypassVal_11 : _GEN_2104; // @[LoadQueue.scala 267:32:@39351.4]
  assign _GEN_2106 = prevPriorityRequest_12 ? io_loadDataFromMem : dataQ_12; // @[LoadQueue.scala 269:44:@39362.6]
  assign _GEN_2107 = bypassRequest_12 ? bypassVal_12 : _GEN_2106; // @[LoadQueue.scala 267:32:@39358.4]
  assign _GEN_2108 = prevPriorityRequest_13 ? io_loadDataFromMem : dataQ_13; // @[LoadQueue.scala 269:44:@39369.6]
  assign _GEN_2109 = bypassRequest_13 ? bypassVal_13 : _GEN_2108; // @[LoadQueue.scala 267:32:@39365.4]
  assign _GEN_2110 = prevPriorityRequest_14 ? io_loadDataFromMem : dataQ_14; // @[LoadQueue.scala 269:44:@39376.6]
  assign _GEN_2111 = bypassRequest_14 ? bypassVal_14 : _GEN_2110; // @[LoadQueue.scala 267:32:@39372.4]
  assign _GEN_2112 = prevPriorityRequest_15 ? io_loadDataFromMem : dataQ_15; // @[LoadQueue.scala 269:44:@39383.6]
  assign _GEN_2113 = bypassRequest_15 ? bypassVal_15 : _GEN_2112; // @[LoadQueue.scala 267:32:@39379.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[LoadQueue.scala 286:69:@39387.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[LoadQueue.scala 286:69:@39389.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[LoadQueue.scala 286:69:@39391.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[LoadQueue.scala 286:69:@39393.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[LoadQueue.scala 286:69:@39395.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[LoadQueue.scala 286:69:@39397.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[LoadQueue.scala 286:69:@39399.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[LoadQueue.scala 286:69:@39401.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[LoadQueue.scala 286:69:@39403.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[LoadQueue.scala 286:69:@39405.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[LoadQueue.scala 286:69:@39407.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[LoadQueue.scala 286:69:@39409.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[LoadQueue.scala 286:69:@39411.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[LoadQueue.scala 286:69:@39413.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[LoadQueue.scala 286:69:@39415.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[LoadQueue.scala 286:69:@39417.4]
  assign _T_94179 = addrKnown_0 == 1'h0; // @[LoadQueue.scala 298:86:@39421.4]
  assign _T_94180 = entriesPorts_0_0 & _T_94179; // @[LoadQueue.scala 298:83:@39422.4]
  assign _T_94182 = addrKnown_1 == 1'h0; // @[LoadQueue.scala 298:86:@39423.4]
  assign _T_94183 = entriesPorts_0_1 & _T_94182; // @[LoadQueue.scala 298:83:@39424.4]
  assign _T_94185 = addrKnown_2 == 1'h0; // @[LoadQueue.scala 298:86:@39425.4]
  assign _T_94186 = entriesPorts_0_2 & _T_94185; // @[LoadQueue.scala 298:83:@39426.4]
  assign _T_94188 = addrKnown_3 == 1'h0; // @[LoadQueue.scala 298:86:@39427.4]
  assign _T_94189 = entriesPorts_0_3 & _T_94188; // @[LoadQueue.scala 298:83:@39428.4]
  assign _T_94191 = addrKnown_4 == 1'h0; // @[LoadQueue.scala 298:86:@39429.4]
  assign _T_94192 = entriesPorts_0_4 & _T_94191; // @[LoadQueue.scala 298:83:@39430.4]
  assign _T_94194 = addrKnown_5 == 1'h0; // @[LoadQueue.scala 298:86:@39431.4]
  assign _T_94195 = entriesPorts_0_5 & _T_94194; // @[LoadQueue.scala 298:83:@39432.4]
  assign _T_94197 = addrKnown_6 == 1'h0; // @[LoadQueue.scala 298:86:@39433.4]
  assign _T_94198 = entriesPorts_0_6 & _T_94197; // @[LoadQueue.scala 298:83:@39434.4]
  assign _T_94200 = addrKnown_7 == 1'h0; // @[LoadQueue.scala 298:86:@39435.4]
  assign _T_94201 = entriesPorts_0_7 & _T_94200; // @[LoadQueue.scala 298:83:@39436.4]
  assign _T_94203 = addrKnown_8 == 1'h0; // @[LoadQueue.scala 298:86:@39437.4]
  assign _T_94204 = entriesPorts_0_8 & _T_94203; // @[LoadQueue.scala 298:83:@39438.4]
  assign _T_94206 = addrKnown_9 == 1'h0; // @[LoadQueue.scala 298:86:@39439.4]
  assign _T_94207 = entriesPorts_0_9 & _T_94206; // @[LoadQueue.scala 298:83:@39440.4]
  assign _T_94209 = addrKnown_10 == 1'h0; // @[LoadQueue.scala 298:86:@39441.4]
  assign _T_94210 = entriesPorts_0_10 & _T_94209; // @[LoadQueue.scala 298:83:@39442.4]
  assign _T_94212 = addrKnown_11 == 1'h0; // @[LoadQueue.scala 298:86:@39443.4]
  assign _T_94213 = entriesPorts_0_11 & _T_94212; // @[LoadQueue.scala 298:83:@39444.4]
  assign _T_94215 = addrKnown_12 == 1'h0; // @[LoadQueue.scala 298:86:@39445.4]
  assign _T_94216 = entriesPorts_0_12 & _T_94215; // @[LoadQueue.scala 298:83:@39446.4]
  assign _T_94218 = addrKnown_13 == 1'h0; // @[LoadQueue.scala 298:86:@39447.4]
  assign _T_94219 = entriesPorts_0_13 & _T_94218; // @[LoadQueue.scala 298:83:@39448.4]
  assign _T_94221 = addrKnown_14 == 1'h0; // @[LoadQueue.scala 298:86:@39449.4]
  assign _T_94222 = entriesPorts_0_14 & _T_94221; // @[LoadQueue.scala 298:83:@39450.4]
  assign _T_94224 = addrKnown_15 == 1'h0; // @[LoadQueue.scala 298:86:@39451.4]
  assign _T_94225 = entriesPorts_0_15 & _T_94224; // @[LoadQueue.scala 298:83:@39452.4]
  assign _T_94308 = _T_94225 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39506.4]
  assign _T_94309 = _T_94222 ? 16'h4000 : _T_94308; // @[Mux.scala 31:69:@39507.4]
  assign _T_94310 = _T_94219 ? 16'h2000 : _T_94309; // @[Mux.scala 31:69:@39508.4]
  assign _T_94311 = _T_94216 ? 16'h1000 : _T_94310; // @[Mux.scala 31:69:@39509.4]
  assign _T_94312 = _T_94213 ? 16'h800 : _T_94311; // @[Mux.scala 31:69:@39510.4]
  assign _T_94313 = _T_94210 ? 16'h400 : _T_94312; // @[Mux.scala 31:69:@39511.4]
  assign _T_94314 = _T_94207 ? 16'h200 : _T_94313; // @[Mux.scala 31:69:@39512.4]
  assign _T_94315 = _T_94204 ? 16'h100 : _T_94314; // @[Mux.scala 31:69:@39513.4]
  assign _T_94316 = _T_94201 ? 16'h80 : _T_94315; // @[Mux.scala 31:69:@39514.4]
  assign _T_94317 = _T_94198 ? 16'h40 : _T_94316; // @[Mux.scala 31:69:@39515.4]
  assign _T_94318 = _T_94195 ? 16'h20 : _T_94317; // @[Mux.scala 31:69:@39516.4]
  assign _T_94319 = _T_94192 ? 16'h10 : _T_94318; // @[Mux.scala 31:69:@39517.4]
  assign _T_94320 = _T_94189 ? 16'h8 : _T_94319; // @[Mux.scala 31:69:@39518.4]
  assign _T_94321 = _T_94186 ? 16'h4 : _T_94320; // @[Mux.scala 31:69:@39519.4]
  assign _T_94322 = _T_94183 ? 16'h2 : _T_94321; // @[Mux.scala 31:69:@39520.4]
  assign _T_94323 = _T_94180 ? 16'h1 : _T_94322; // @[Mux.scala 31:69:@39521.4]
  assign _T_94324 = _T_94323[0]; // @[OneHot.scala 66:30:@39522.4]
  assign _T_94325 = _T_94323[1]; // @[OneHot.scala 66:30:@39523.4]
  assign _T_94326 = _T_94323[2]; // @[OneHot.scala 66:30:@39524.4]
  assign _T_94327 = _T_94323[3]; // @[OneHot.scala 66:30:@39525.4]
  assign _T_94328 = _T_94323[4]; // @[OneHot.scala 66:30:@39526.4]
  assign _T_94329 = _T_94323[5]; // @[OneHot.scala 66:30:@39527.4]
  assign _T_94330 = _T_94323[6]; // @[OneHot.scala 66:30:@39528.4]
  assign _T_94331 = _T_94323[7]; // @[OneHot.scala 66:30:@39529.4]
  assign _T_94332 = _T_94323[8]; // @[OneHot.scala 66:30:@39530.4]
  assign _T_94333 = _T_94323[9]; // @[OneHot.scala 66:30:@39531.4]
  assign _T_94334 = _T_94323[10]; // @[OneHot.scala 66:30:@39532.4]
  assign _T_94335 = _T_94323[11]; // @[OneHot.scala 66:30:@39533.4]
  assign _T_94336 = _T_94323[12]; // @[OneHot.scala 66:30:@39534.4]
  assign _T_94337 = _T_94323[13]; // @[OneHot.scala 66:30:@39535.4]
  assign _T_94338 = _T_94323[14]; // @[OneHot.scala 66:30:@39536.4]
  assign _T_94339 = _T_94323[15]; // @[OneHot.scala 66:30:@39537.4]
  assign _T_94380 = _T_94180 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39555.4]
  assign _T_94381 = _T_94225 ? 16'h4000 : _T_94380; // @[Mux.scala 31:69:@39556.4]
  assign _T_94382 = _T_94222 ? 16'h2000 : _T_94381; // @[Mux.scala 31:69:@39557.4]
  assign _T_94383 = _T_94219 ? 16'h1000 : _T_94382; // @[Mux.scala 31:69:@39558.4]
  assign _T_94384 = _T_94216 ? 16'h800 : _T_94383; // @[Mux.scala 31:69:@39559.4]
  assign _T_94385 = _T_94213 ? 16'h400 : _T_94384; // @[Mux.scala 31:69:@39560.4]
  assign _T_94386 = _T_94210 ? 16'h200 : _T_94385; // @[Mux.scala 31:69:@39561.4]
  assign _T_94387 = _T_94207 ? 16'h100 : _T_94386; // @[Mux.scala 31:69:@39562.4]
  assign _T_94388 = _T_94204 ? 16'h80 : _T_94387; // @[Mux.scala 31:69:@39563.4]
  assign _T_94389 = _T_94201 ? 16'h40 : _T_94388; // @[Mux.scala 31:69:@39564.4]
  assign _T_94390 = _T_94198 ? 16'h20 : _T_94389; // @[Mux.scala 31:69:@39565.4]
  assign _T_94391 = _T_94195 ? 16'h10 : _T_94390; // @[Mux.scala 31:69:@39566.4]
  assign _T_94392 = _T_94192 ? 16'h8 : _T_94391; // @[Mux.scala 31:69:@39567.4]
  assign _T_94393 = _T_94189 ? 16'h4 : _T_94392; // @[Mux.scala 31:69:@39568.4]
  assign _T_94394 = _T_94186 ? 16'h2 : _T_94393; // @[Mux.scala 31:69:@39569.4]
  assign _T_94395 = _T_94183 ? 16'h1 : _T_94394; // @[Mux.scala 31:69:@39570.4]
  assign _T_94396 = _T_94395[0]; // @[OneHot.scala 66:30:@39571.4]
  assign _T_94397 = _T_94395[1]; // @[OneHot.scala 66:30:@39572.4]
  assign _T_94398 = _T_94395[2]; // @[OneHot.scala 66:30:@39573.4]
  assign _T_94399 = _T_94395[3]; // @[OneHot.scala 66:30:@39574.4]
  assign _T_94400 = _T_94395[4]; // @[OneHot.scala 66:30:@39575.4]
  assign _T_94401 = _T_94395[5]; // @[OneHot.scala 66:30:@39576.4]
  assign _T_94402 = _T_94395[6]; // @[OneHot.scala 66:30:@39577.4]
  assign _T_94403 = _T_94395[7]; // @[OneHot.scala 66:30:@39578.4]
  assign _T_94404 = _T_94395[8]; // @[OneHot.scala 66:30:@39579.4]
  assign _T_94405 = _T_94395[9]; // @[OneHot.scala 66:30:@39580.4]
  assign _T_94406 = _T_94395[10]; // @[OneHot.scala 66:30:@39581.4]
  assign _T_94407 = _T_94395[11]; // @[OneHot.scala 66:30:@39582.4]
  assign _T_94408 = _T_94395[12]; // @[OneHot.scala 66:30:@39583.4]
  assign _T_94409 = _T_94395[13]; // @[OneHot.scala 66:30:@39584.4]
  assign _T_94410 = _T_94395[14]; // @[OneHot.scala 66:30:@39585.4]
  assign _T_94411 = _T_94395[15]; // @[OneHot.scala 66:30:@39586.4]
  assign _T_94452 = _T_94183 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39604.4]
  assign _T_94453 = _T_94180 ? 16'h4000 : _T_94452; // @[Mux.scala 31:69:@39605.4]
  assign _T_94454 = _T_94225 ? 16'h2000 : _T_94453; // @[Mux.scala 31:69:@39606.4]
  assign _T_94455 = _T_94222 ? 16'h1000 : _T_94454; // @[Mux.scala 31:69:@39607.4]
  assign _T_94456 = _T_94219 ? 16'h800 : _T_94455; // @[Mux.scala 31:69:@39608.4]
  assign _T_94457 = _T_94216 ? 16'h400 : _T_94456; // @[Mux.scala 31:69:@39609.4]
  assign _T_94458 = _T_94213 ? 16'h200 : _T_94457; // @[Mux.scala 31:69:@39610.4]
  assign _T_94459 = _T_94210 ? 16'h100 : _T_94458; // @[Mux.scala 31:69:@39611.4]
  assign _T_94460 = _T_94207 ? 16'h80 : _T_94459; // @[Mux.scala 31:69:@39612.4]
  assign _T_94461 = _T_94204 ? 16'h40 : _T_94460; // @[Mux.scala 31:69:@39613.4]
  assign _T_94462 = _T_94201 ? 16'h20 : _T_94461; // @[Mux.scala 31:69:@39614.4]
  assign _T_94463 = _T_94198 ? 16'h10 : _T_94462; // @[Mux.scala 31:69:@39615.4]
  assign _T_94464 = _T_94195 ? 16'h8 : _T_94463; // @[Mux.scala 31:69:@39616.4]
  assign _T_94465 = _T_94192 ? 16'h4 : _T_94464; // @[Mux.scala 31:69:@39617.4]
  assign _T_94466 = _T_94189 ? 16'h2 : _T_94465; // @[Mux.scala 31:69:@39618.4]
  assign _T_94467 = _T_94186 ? 16'h1 : _T_94466; // @[Mux.scala 31:69:@39619.4]
  assign _T_94468 = _T_94467[0]; // @[OneHot.scala 66:30:@39620.4]
  assign _T_94469 = _T_94467[1]; // @[OneHot.scala 66:30:@39621.4]
  assign _T_94470 = _T_94467[2]; // @[OneHot.scala 66:30:@39622.4]
  assign _T_94471 = _T_94467[3]; // @[OneHot.scala 66:30:@39623.4]
  assign _T_94472 = _T_94467[4]; // @[OneHot.scala 66:30:@39624.4]
  assign _T_94473 = _T_94467[5]; // @[OneHot.scala 66:30:@39625.4]
  assign _T_94474 = _T_94467[6]; // @[OneHot.scala 66:30:@39626.4]
  assign _T_94475 = _T_94467[7]; // @[OneHot.scala 66:30:@39627.4]
  assign _T_94476 = _T_94467[8]; // @[OneHot.scala 66:30:@39628.4]
  assign _T_94477 = _T_94467[9]; // @[OneHot.scala 66:30:@39629.4]
  assign _T_94478 = _T_94467[10]; // @[OneHot.scala 66:30:@39630.4]
  assign _T_94479 = _T_94467[11]; // @[OneHot.scala 66:30:@39631.4]
  assign _T_94480 = _T_94467[12]; // @[OneHot.scala 66:30:@39632.4]
  assign _T_94481 = _T_94467[13]; // @[OneHot.scala 66:30:@39633.4]
  assign _T_94482 = _T_94467[14]; // @[OneHot.scala 66:30:@39634.4]
  assign _T_94483 = _T_94467[15]; // @[OneHot.scala 66:30:@39635.4]
  assign _T_94524 = _T_94186 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39653.4]
  assign _T_94525 = _T_94183 ? 16'h4000 : _T_94524; // @[Mux.scala 31:69:@39654.4]
  assign _T_94526 = _T_94180 ? 16'h2000 : _T_94525; // @[Mux.scala 31:69:@39655.4]
  assign _T_94527 = _T_94225 ? 16'h1000 : _T_94526; // @[Mux.scala 31:69:@39656.4]
  assign _T_94528 = _T_94222 ? 16'h800 : _T_94527; // @[Mux.scala 31:69:@39657.4]
  assign _T_94529 = _T_94219 ? 16'h400 : _T_94528; // @[Mux.scala 31:69:@39658.4]
  assign _T_94530 = _T_94216 ? 16'h200 : _T_94529; // @[Mux.scala 31:69:@39659.4]
  assign _T_94531 = _T_94213 ? 16'h100 : _T_94530; // @[Mux.scala 31:69:@39660.4]
  assign _T_94532 = _T_94210 ? 16'h80 : _T_94531; // @[Mux.scala 31:69:@39661.4]
  assign _T_94533 = _T_94207 ? 16'h40 : _T_94532; // @[Mux.scala 31:69:@39662.4]
  assign _T_94534 = _T_94204 ? 16'h20 : _T_94533; // @[Mux.scala 31:69:@39663.4]
  assign _T_94535 = _T_94201 ? 16'h10 : _T_94534; // @[Mux.scala 31:69:@39664.4]
  assign _T_94536 = _T_94198 ? 16'h8 : _T_94535; // @[Mux.scala 31:69:@39665.4]
  assign _T_94537 = _T_94195 ? 16'h4 : _T_94536; // @[Mux.scala 31:69:@39666.4]
  assign _T_94538 = _T_94192 ? 16'h2 : _T_94537; // @[Mux.scala 31:69:@39667.4]
  assign _T_94539 = _T_94189 ? 16'h1 : _T_94538; // @[Mux.scala 31:69:@39668.4]
  assign _T_94540 = _T_94539[0]; // @[OneHot.scala 66:30:@39669.4]
  assign _T_94541 = _T_94539[1]; // @[OneHot.scala 66:30:@39670.4]
  assign _T_94542 = _T_94539[2]; // @[OneHot.scala 66:30:@39671.4]
  assign _T_94543 = _T_94539[3]; // @[OneHot.scala 66:30:@39672.4]
  assign _T_94544 = _T_94539[4]; // @[OneHot.scala 66:30:@39673.4]
  assign _T_94545 = _T_94539[5]; // @[OneHot.scala 66:30:@39674.4]
  assign _T_94546 = _T_94539[6]; // @[OneHot.scala 66:30:@39675.4]
  assign _T_94547 = _T_94539[7]; // @[OneHot.scala 66:30:@39676.4]
  assign _T_94548 = _T_94539[8]; // @[OneHot.scala 66:30:@39677.4]
  assign _T_94549 = _T_94539[9]; // @[OneHot.scala 66:30:@39678.4]
  assign _T_94550 = _T_94539[10]; // @[OneHot.scala 66:30:@39679.4]
  assign _T_94551 = _T_94539[11]; // @[OneHot.scala 66:30:@39680.4]
  assign _T_94552 = _T_94539[12]; // @[OneHot.scala 66:30:@39681.4]
  assign _T_94553 = _T_94539[13]; // @[OneHot.scala 66:30:@39682.4]
  assign _T_94554 = _T_94539[14]; // @[OneHot.scala 66:30:@39683.4]
  assign _T_94555 = _T_94539[15]; // @[OneHot.scala 66:30:@39684.4]
  assign _T_94596 = _T_94189 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39702.4]
  assign _T_94597 = _T_94186 ? 16'h4000 : _T_94596; // @[Mux.scala 31:69:@39703.4]
  assign _T_94598 = _T_94183 ? 16'h2000 : _T_94597; // @[Mux.scala 31:69:@39704.4]
  assign _T_94599 = _T_94180 ? 16'h1000 : _T_94598; // @[Mux.scala 31:69:@39705.4]
  assign _T_94600 = _T_94225 ? 16'h800 : _T_94599; // @[Mux.scala 31:69:@39706.4]
  assign _T_94601 = _T_94222 ? 16'h400 : _T_94600; // @[Mux.scala 31:69:@39707.4]
  assign _T_94602 = _T_94219 ? 16'h200 : _T_94601; // @[Mux.scala 31:69:@39708.4]
  assign _T_94603 = _T_94216 ? 16'h100 : _T_94602; // @[Mux.scala 31:69:@39709.4]
  assign _T_94604 = _T_94213 ? 16'h80 : _T_94603; // @[Mux.scala 31:69:@39710.4]
  assign _T_94605 = _T_94210 ? 16'h40 : _T_94604; // @[Mux.scala 31:69:@39711.4]
  assign _T_94606 = _T_94207 ? 16'h20 : _T_94605; // @[Mux.scala 31:69:@39712.4]
  assign _T_94607 = _T_94204 ? 16'h10 : _T_94606; // @[Mux.scala 31:69:@39713.4]
  assign _T_94608 = _T_94201 ? 16'h8 : _T_94607; // @[Mux.scala 31:69:@39714.4]
  assign _T_94609 = _T_94198 ? 16'h4 : _T_94608; // @[Mux.scala 31:69:@39715.4]
  assign _T_94610 = _T_94195 ? 16'h2 : _T_94609; // @[Mux.scala 31:69:@39716.4]
  assign _T_94611 = _T_94192 ? 16'h1 : _T_94610; // @[Mux.scala 31:69:@39717.4]
  assign _T_94612 = _T_94611[0]; // @[OneHot.scala 66:30:@39718.4]
  assign _T_94613 = _T_94611[1]; // @[OneHot.scala 66:30:@39719.4]
  assign _T_94614 = _T_94611[2]; // @[OneHot.scala 66:30:@39720.4]
  assign _T_94615 = _T_94611[3]; // @[OneHot.scala 66:30:@39721.4]
  assign _T_94616 = _T_94611[4]; // @[OneHot.scala 66:30:@39722.4]
  assign _T_94617 = _T_94611[5]; // @[OneHot.scala 66:30:@39723.4]
  assign _T_94618 = _T_94611[6]; // @[OneHot.scala 66:30:@39724.4]
  assign _T_94619 = _T_94611[7]; // @[OneHot.scala 66:30:@39725.4]
  assign _T_94620 = _T_94611[8]; // @[OneHot.scala 66:30:@39726.4]
  assign _T_94621 = _T_94611[9]; // @[OneHot.scala 66:30:@39727.4]
  assign _T_94622 = _T_94611[10]; // @[OneHot.scala 66:30:@39728.4]
  assign _T_94623 = _T_94611[11]; // @[OneHot.scala 66:30:@39729.4]
  assign _T_94624 = _T_94611[12]; // @[OneHot.scala 66:30:@39730.4]
  assign _T_94625 = _T_94611[13]; // @[OneHot.scala 66:30:@39731.4]
  assign _T_94626 = _T_94611[14]; // @[OneHot.scala 66:30:@39732.4]
  assign _T_94627 = _T_94611[15]; // @[OneHot.scala 66:30:@39733.4]
  assign _T_94668 = _T_94192 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39751.4]
  assign _T_94669 = _T_94189 ? 16'h4000 : _T_94668; // @[Mux.scala 31:69:@39752.4]
  assign _T_94670 = _T_94186 ? 16'h2000 : _T_94669; // @[Mux.scala 31:69:@39753.4]
  assign _T_94671 = _T_94183 ? 16'h1000 : _T_94670; // @[Mux.scala 31:69:@39754.4]
  assign _T_94672 = _T_94180 ? 16'h800 : _T_94671; // @[Mux.scala 31:69:@39755.4]
  assign _T_94673 = _T_94225 ? 16'h400 : _T_94672; // @[Mux.scala 31:69:@39756.4]
  assign _T_94674 = _T_94222 ? 16'h200 : _T_94673; // @[Mux.scala 31:69:@39757.4]
  assign _T_94675 = _T_94219 ? 16'h100 : _T_94674; // @[Mux.scala 31:69:@39758.4]
  assign _T_94676 = _T_94216 ? 16'h80 : _T_94675; // @[Mux.scala 31:69:@39759.4]
  assign _T_94677 = _T_94213 ? 16'h40 : _T_94676; // @[Mux.scala 31:69:@39760.4]
  assign _T_94678 = _T_94210 ? 16'h20 : _T_94677; // @[Mux.scala 31:69:@39761.4]
  assign _T_94679 = _T_94207 ? 16'h10 : _T_94678; // @[Mux.scala 31:69:@39762.4]
  assign _T_94680 = _T_94204 ? 16'h8 : _T_94679; // @[Mux.scala 31:69:@39763.4]
  assign _T_94681 = _T_94201 ? 16'h4 : _T_94680; // @[Mux.scala 31:69:@39764.4]
  assign _T_94682 = _T_94198 ? 16'h2 : _T_94681; // @[Mux.scala 31:69:@39765.4]
  assign _T_94683 = _T_94195 ? 16'h1 : _T_94682; // @[Mux.scala 31:69:@39766.4]
  assign _T_94684 = _T_94683[0]; // @[OneHot.scala 66:30:@39767.4]
  assign _T_94685 = _T_94683[1]; // @[OneHot.scala 66:30:@39768.4]
  assign _T_94686 = _T_94683[2]; // @[OneHot.scala 66:30:@39769.4]
  assign _T_94687 = _T_94683[3]; // @[OneHot.scala 66:30:@39770.4]
  assign _T_94688 = _T_94683[4]; // @[OneHot.scala 66:30:@39771.4]
  assign _T_94689 = _T_94683[5]; // @[OneHot.scala 66:30:@39772.4]
  assign _T_94690 = _T_94683[6]; // @[OneHot.scala 66:30:@39773.4]
  assign _T_94691 = _T_94683[7]; // @[OneHot.scala 66:30:@39774.4]
  assign _T_94692 = _T_94683[8]; // @[OneHot.scala 66:30:@39775.4]
  assign _T_94693 = _T_94683[9]; // @[OneHot.scala 66:30:@39776.4]
  assign _T_94694 = _T_94683[10]; // @[OneHot.scala 66:30:@39777.4]
  assign _T_94695 = _T_94683[11]; // @[OneHot.scala 66:30:@39778.4]
  assign _T_94696 = _T_94683[12]; // @[OneHot.scala 66:30:@39779.4]
  assign _T_94697 = _T_94683[13]; // @[OneHot.scala 66:30:@39780.4]
  assign _T_94698 = _T_94683[14]; // @[OneHot.scala 66:30:@39781.4]
  assign _T_94699 = _T_94683[15]; // @[OneHot.scala 66:30:@39782.4]
  assign _T_94740 = _T_94195 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39800.4]
  assign _T_94741 = _T_94192 ? 16'h4000 : _T_94740; // @[Mux.scala 31:69:@39801.4]
  assign _T_94742 = _T_94189 ? 16'h2000 : _T_94741; // @[Mux.scala 31:69:@39802.4]
  assign _T_94743 = _T_94186 ? 16'h1000 : _T_94742; // @[Mux.scala 31:69:@39803.4]
  assign _T_94744 = _T_94183 ? 16'h800 : _T_94743; // @[Mux.scala 31:69:@39804.4]
  assign _T_94745 = _T_94180 ? 16'h400 : _T_94744; // @[Mux.scala 31:69:@39805.4]
  assign _T_94746 = _T_94225 ? 16'h200 : _T_94745; // @[Mux.scala 31:69:@39806.4]
  assign _T_94747 = _T_94222 ? 16'h100 : _T_94746; // @[Mux.scala 31:69:@39807.4]
  assign _T_94748 = _T_94219 ? 16'h80 : _T_94747; // @[Mux.scala 31:69:@39808.4]
  assign _T_94749 = _T_94216 ? 16'h40 : _T_94748; // @[Mux.scala 31:69:@39809.4]
  assign _T_94750 = _T_94213 ? 16'h20 : _T_94749; // @[Mux.scala 31:69:@39810.4]
  assign _T_94751 = _T_94210 ? 16'h10 : _T_94750; // @[Mux.scala 31:69:@39811.4]
  assign _T_94752 = _T_94207 ? 16'h8 : _T_94751; // @[Mux.scala 31:69:@39812.4]
  assign _T_94753 = _T_94204 ? 16'h4 : _T_94752; // @[Mux.scala 31:69:@39813.4]
  assign _T_94754 = _T_94201 ? 16'h2 : _T_94753; // @[Mux.scala 31:69:@39814.4]
  assign _T_94755 = _T_94198 ? 16'h1 : _T_94754; // @[Mux.scala 31:69:@39815.4]
  assign _T_94756 = _T_94755[0]; // @[OneHot.scala 66:30:@39816.4]
  assign _T_94757 = _T_94755[1]; // @[OneHot.scala 66:30:@39817.4]
  assign _T_94758 = _T_94755[2]; // @[OneHot.scala 66:30:@39818.4]
  assign _T_94759 = _T_94755[3]; // @[OneHot.scala 66:30:@39819.4]
  assign _T_94760 = _T_94755[4]; // @[OneHot.scala 66:30:@39820.4]
  assign _T_94761 = _T_94755[5]; // @[OneHot.scala 66:30:@39821.4]
  assign _T_94762 = _T_94755[6]; // @[OneHot.scala 66:30:@39822.4]
  assign _T_94763 = _T_94755[7]; // @[OneHot.scala 66:30:@39823.4]
  assign _T_94764 = _T_94755[8]; // @[OneHot.scala 66:30:@39824.4]
  assign _T_94765 = _T_94755[9]; // @[OneHot.scala 66:30:@39825.4]
  assign _T_94766 = _T_94755[10]; // @[OneHot.scala 66:30:@39826.4]
  assign _T_94767 = _T_94755[11]; // @[OneHot.scala 66:30:@39827.4]
  assign _T_94768 = _T_94755[12]; // @[OneHot.scala 66:30:@39828.4]
  assign _T_94769 = _T_94755[13]; // @[OneHot.scala 66:30:@39829.4]
  assign _T_94770 = _T_94755[14]; // @[OneHot.scala 66:30:@39830.4]
  assign _T_94771 = _T_94755[15]; // @[OneHot.scala 66:30:@39831.4]
  assign _T_94812 = _T_94198 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39849.4]
  assign _T_94813 = _T_94195 ? 16'h4000 : _T_94812; // @[Mux.scala 31:69:@39850.4]
  assign _T_94814 = _T_94192 ? 16'h2000 : _T_94813; // @[Mux.scala 31:69:@39851.4]
  assign _T_94815 = _T_94189 ? 16'h1000 : _T_94814; // @[Mux.scala 31:69:@39852.4]
  assign _T_94816 = _T_94186 ? 16'h800 : _T_94815; // @[Mux.scala 31:69:@39853.4]
  assign _T_94817 = _T_94183 ? 16'h400 : _T_94816; // @[Mux.scala 31:69:@39854.4]
  assign _T_94818 = _T_94180 ? 16'h200 : _T_94817; // @[Mux.scala 31:69:@39855.4]
  assign _T_94819 = _T_94225 ? 16'h100 : _T_94818; // @[Mux.scala 31:69:@39856.4]
  assign _T_94820 = _T_94222 ? 16'h80 : _T_94819; // @[Mux.scala 31:69:@39857.4]
  assign _T_94821 = _T_94219 ? 16'h40 : _T_94820; // @[Mux.scala 31:69:@39858.4]
  assign _T_94822 = _T_94216 ? 16'h20 : _T_94821; // @[Mux.scala 31:69:@39859.4]
  assign _T_94823 = _T_94213 ? 16'h10 : _T_94822; // @[Mux.scala 31:69:@39860.4]
  assign _T_94824 = _T_94210 ? 16'h8 : _T_94823; // @[Mux.scala 31:69:@39861.4]
  assign _T_94825 = _T_94207 ? 16'h4 : _T_94824; // @[Mux.scala 31:69:@39862.4]
  assign _T_94826 = _T_94204 ? 16'h2 : _T_94825; // @[Mux.scala 31:69:@39863.4]
  assign _T_94827 = _T_94201 ? 16'h1 : _T_94826; // @[Mux.scala 31:69:@39864.4]
  assign _T_94828 = _T_94827[0]; // @[OneHot.scala 66:30:@39865.4]
  assign _T_94829 = _T_94827[1]; // @[OneHot.scala 66:30:@39866.4]
  assign _T_94830 = _T_94827[2]; // @[OneHot.scala 66:30:@39867.4]
  assign _T_94831 = _T_94827[3]; // @[OneHot.scala 66:30:@39868.4]
  assign _T_94832 = _T_94827[4]; // @[OneHot.scala 66:30:@39869.4]
  assign _T_94833 = _T_94827[5]; // @[OneHot.scala 66:30:@39870.4]
  assign _T_94834 = _T_94827[6]; // @[OneHot.scala 66:30:@39871.4]
  assign _T_94835 = _T_94827[7]; // @[OneHot.scala 66:30:@39872.4]
  assign _T_94836 = _T_94827[8]; // @[OneHot.scala 66:30:@39873.4]
  assign _T_94837 = _T_94827[9]; // @[OneHot.scala 66:30:@39874.4]
  assign _T_94838 = _T_94827[10]; // @[OneHot.scala 66:30:@39875.4]
  assign _T_94839 = _T_94827[11]; // @[OneHot.scala 66:30:@39876.4]
  assign _T_94840 = _T_94827[12]; // @[OneHot.scala 66:30:@39877.4]
  assign _T_94841 = _T_94827[13]; // @[OneHot.scala 66:30:@39878.4]
  assign _T_94842 = _T_94827[14]; // @[OneHot.scala 66:30:@39879.4]
  assign _T_94843 = _T_94827[15]; // @[OneHot.scala 66:30:@39880.4]
  assign _T_94884 = _T_94201 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39898.4]
  assign _T_94885 = _T_94198 ? 16'h4000 : _T_94884; // @[Mux.scala 31:69:@39899.4]
  assign _T_94886 = _T_94195 ? 16'h2000 : _T_94885; // @[Mux.scala 31:69:@39900.4]
  assign _T_94887 = _T_94192 ? 16'h1000 : _T_94886; // @[Mux.scala 31:69:@39901.4]
  assign _T_94888 = _T_94189 ? 16'h800 : _T_94887; // @[Mux.scala 31:69:@39902.4]
  assign _T_94889 = _T_94186 ? 16'h400 : _T_94888; // @[Mux.scala 31:69:@39903.4]
  assign _T_94890 = _T_94183 ? 16'h200 : _T_94889; // @[Mux.scala 31:69:@39904.4]
  assign _T_94891 = _T_94180 ? 16'h100 : _T_94890; // @[Mux.scala 31:69:@39905.4]
  assign _T_94892 = _T_94225 ? 16'h80 : _T_94891; // @[Mux.scala 31:69:@39906.4]
  assign _T_94893 = _T_94222 ? 16'h40 : _T_94892; // @[Mux.scala 31:69:@39907.4]
  assign _T_94894 = _T_94219 ? 16'h20 : _T_94893; // @[Mux.scala 31:69:@39908.4]
  assign _T_94895 = _T_94216 ? 16'h10 : _T_94894; // @[Mux.scala 31:69:@39909.4]
  assign _T_94896 = _T_94213 ? 16'h8 : _T_94895; // @[Mux.scala 31:69:@39910.4]
  assign _T_94897 = _T_94210 ? 16'h4 : _T_94896; // @[Mux.scala 31:69:@39911.4]
  assign _T_94898 = _T_94207 ? 16'h2 : _T_94897; // @[Mux.scala 31:69:@39912.4]
  assign _T_94899 = _T_94204 ? 16'h1 : _T_94898; // @[Mux.scala 31:69:@39913.4]
  assign _T_94900 = _T_94899[0]; // @[OneHot.scala 66:30:@39914.4]
  assign _T_94901 = _T_94899[1]; // @[OneHot.scala 66:30:@39915.4]
  assign _T_94902 = _T_94899[2]; // @[OneHot.scala 66:30:@39916.4]
  assign _T_94903 = _T_94899[3]; // @[OneHot.scala 66:30:@39917.4]
  assign _T_94904 = _T_94899[4]; // @[OneHot.scala 66:30:@39918.4]
  assign _T_94905 = _T_94899[5]; // @[OneHot.scala 66:30:@39919.4]
  assign _T_94906 = _T_94899[6]; // @[OneHot.scala 66:30:@39920.4]
  assign _T_94907 = _T_94899[7]; // @[OneHot.scala 66:30:@39921.4]
  assign _T_94908 = _T_94899[8]; // @[OneHot.scala 66:30:@39922.4]
  assign _T_94909 = _T_94899[9]; // @[OneHot.scala 66:30:@39923.4]
  assign _T_94910 = _T_94899[10]; // @[OneHot.scala 66:30:@39924.4]
  assign _T_94911 = _T_94899[11]; // @[OneHot.scala 66:30:@39925.4]
  assign _T_94912 = _T_94899[12]; // @[OneHot.scala 66:30:@39926.4]
  assign _T_94913 = _T_94899[13]; // @[OneHot.scala 66:30:@39927.4]
  assign _T_94914 = _T_94899[14]; // @[OneHot.scala 66:30:@39928.4]
  assign _T_94915 = _T_94899[15]; // @[OneHot.scala 66:30:@39929.4]
  assign _T_94956 = _T_94204 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39947.4]
  assign _T_94957 = _T_94201 ? 16'h4000 : _T_94956; // @[Mux.scala 31:69:@39948.4]
  assign _T_94958 = _T_94198 ? 16'h2000 : _T_94957; // @[Mux.scala 31:69:@39949.4]
  assign _T_94959 = _T_94195 ? 16'h1000 : _T_94958; // @[Mux.scala 31:69:@39950.4]
  assign _T_94960 = _T_94192 ? 16'h800 : _T_94959; // @[Mux.scala 31:69:@39951.4]
  assign _T_94961 = _T_94189 ? 16'h400 : _T_94960; // @[Mux.scala 31:69:@39952.4]
  assign _T_94962 = _T_94186 ? 16'h200 : _T_94961; // @[Mux.scala 31:69:@39953.4]
  assign _T_94963 = _T_94183 ? 16'h100 : _T_94962; // @[Mux.scala 31:69:@39954.4]
  assign _T_94964 = _T_94180 ? 16'h80 : _T_94963; // @[Mux.scala 31:69:@39955.4]
  assign _T_94965 = _T_94225 ? 16'h40 : _T_94964; // @[Mux.scala 31:69:@39956.4]
  assign _T_94966 = _T_94222 ? 16'h20 : _T_94965; // @[Mux.scala 31:69:@39957.4]
  assign _T_94967 = _T_94219 ? 16'h10 : _T_94966; // @[Mux.scala 31:69:@39958.4]
  assign _T_94968 = _T_94216 ? 16'h8 : _T_94967; // @[Mux.scala 31:69:@39959.4]
  assign _T_94969 = _T_94213 ? 16'h4 : _T_94968; // @[Mux.scala 31:69:@39960.4]
  assign _T_94970 = _T_94210 ? 16'h2 : _T_94969; // @[Mux.scala 31:69:@39961.4]
  assign _T_94971 = _T_94207 ? 16'h1 : _T_94970; // @[Mux.scala 31:69:@39962.4]
  assign _T_94972 = _T_94971[0]; // @[OneHot.scala 66:30:@39963.4]
  assign _T_94973 = _T_94971[1]; // @[OneHot.scala 66:30:@39964.4]
  assign _T_94974 = _T_94971[2]; // @[OneHot.scala 66:30:@39965.4]
  assign _T_94975 = _T_94971[3]; // @[OneHot.scala 66:30:@39966.4]
  assign _T_94976 = _T_94971[4]; // @[OneHot.scala 66:30:@39967.4]
  assign _T_94977 = _T_94971[5]; // @[OneHot.scala 66:30:@39968.4]
  assign _T_94978 = _T_94971[6]; // @[OneHot.scala 66:30:@39969.4]
  assign _T_94979 = _T_94971[7]; // @[OneHot.scala 66:30:@39970.4]
  assign _T_94980 = _T_94971[8]; // @[OneHot.scala 66:30:@39971.4]
  assign _T_94981 = _T_94971[9]; // @[OneHot.scala 66:30:@39972.4]
  assign _T_94982 = _T_94971[10]; // @[OneHot.scala 66:30:@39973.4]
  assign _T_94983 = _T_94971[11]; // @[OneHot.scala 66:30:@39974.4]
  assign _T_94984 = _T_94971[12]; // @[OneHot.scala 66:30:@39975.4]
  assign _T_94985 = _T_94971[13]; // @[OneHot.scala 66:30:@39976.4]
  assign _T_94986 = _T_94971[14]; // @[OneHot.scala 66:30:@39977.4]
  assign _T_94987 = _T_94971[15]; // @[OneHot.scala 66:30:@39978.4]
  assign _T_95028 = _T_94207 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39996.4]
  assign _T_95029 = _T_94204 ? 16'h4000 : _T_95028; // @[Mux.scala 31:69:@39997.4]
  assign _T_95030 = _T_94201 ? 16'h2000 : _T_95029; // @[Mux.scala 31:69:@39998.4]
  assign _T_95031 = _T_94198 ? 16'h1000 : _T_95030; // @[Mux.scala 31:69:@39999.4]
  assign _T_95032 = _T_94195 ? 16'h800 : _T_95031; // @[Mux.scala 31:69:@40000.4]
  assign _T_95033 = _T_94192 ? 16'h400 : _T_95032; // @[Mux.scala 31:69:@40001.4]
  assign _T_95034 = _T_94189 ? 16'h200 : _T_95033; // @[Mux.scala 31:69:@40002.4]
  assign _T_95035 = _T_94186 ? 16'h100 : _T_95034; // @[Mux.scala 31:69:@40003.4]
  assign _T_95036 = _T_94183 ? 16'h80 : _T_95035; // @[Mux.scala 31:69:@40004.4]
  assign _T_95037 = _T_94180 ? 16'h40 : _T_95036; // @[Mux.scala 31:69:@40005.4]
  assign _T_95038 = _T_94225 ? 16'h20 : _T_95037; // @[Mux.scala 31:69:@40006.4]
  assign _T_95039 = _T_94222 ? 16'h10 : _T_95038; // @[Mux.scala 31:69:@40007.4]
  assign _T_95040 = _T_94219 ? 16'h8 : _T_95039; // @[Mux.scala 31:69:@40008.4]
  assign _T_95041 = _T_94216 ? 16'h4 : _T_95040; // @[Mux.scala 31:69:@40009.4]
  assign _T_95042 = _T_94213 ? 16'h2 : _T_95041; // @[Mux.scala 31:69:@40010.4]
  assign _T_95043 = _T_94210 ? 16'h1 : _T_95042; // @[Mux.scala 31:69:@40011.4]
  assign _T_95044 = _T_95043[0]; // @[OneHot.scala 66:30:@40012.4]
  assign _T_95045 = _T_95043[1]; // @[OneHot.scala 66:30:@40013.4]
  assign _T_95046 = _T_95043[2]; // @[OneHot.scala 66:30:@40014.4]
  assign _T_95047 = _T_95043[3]; // @[OneHot.scala 66:30:@40015.4]
  assign _T_95048 = _T_95043[4]; // @[OneHot.scala 66:30:@40016.4]
  assign _T_95049 = _T_95043[5]; // @[OneHot.scala 66:30:@40017.4]
  assign _T_95050 = _T_95043[6]; // @[OneHot.scala 66:30:@40018.4]
  assign _T_95051 = _T_95043[7]; // @[OneHot.scala 66:30:@40019.4]
  assign _T_95052 = _T_95043[8]; // @[OneHot.scala 66:30:@40020.4]
  assign _T_95053 = _T_95043[9]; // @[OneHot.scala 66:30:@40021.4]
  assign _T_95054 = _T_95043[10]; // @[OneHot.scala 66:30:@40022.4]
  assign _T_95055 = _T_95043[11]; // @[OneHot.scala 66:30:@40023.4]
  assign _T_95056 = _T_95043[12]; // @[OneHot.scala 66:30:@40024.4]
  assign _T_95057 = _T_95043[13]; // @[OneHot.scala 66:30:@40025.4]
  assign _T_95058 = _T_95043[14]; // @[OneHot.scala 66:30:@40026.4]
  assign _T_95059 = _T_95043[15]; // @[OneHot.scala 66:30:@40027.4]
  assign _T_95100 = _T_94210 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40045.4]
  assign _T_95101 = _T_94207 ? 16'h4000 : _T_95100; // @[Mux.scala 31:69:@40046.4]
  assign _T_95102 = _T_94204 ? 16'h2000 : _T_95101; // @[Mux.scala 31:69:@40047.4]
  assign _T_95103 = _T_94201 ? 16'h1000 : _T_95102; // @[Mux.scala 31:69:@40048.4]
  assign _T_95104 = _T_94198 ? 16'h800 : _T_95103; // @[Mux.scala 31:69:@40049.4]
  assign _T_95105 = _T_94195 ? 16'h400 : _T_95104; // @[Mux.scala 31:69:@40050.4]
  assign _T_95106 = _T_94192 ? 16'h200 : _T_95105; // @[Mux.scala 31:69:@40051.4]
  assign _T_95107 = _T_94189 ? 16'h100 : _T_95106; // @[Mux.scala 31:69:@40052.4]
  assign _T_95108 = _T_94186 ? 16'h80 : _T_95107; // @[Mux.scala 31:69:@40053.4]
  assign _T_95109 = _T_94183 ? 16'h40 : _T_95108; // @[Mux.scala 31:69:@40054.4]
  assign _T_95110 = _T_94180 ? 16'h20 : _T_95109; // @[Mux.scala 31:69:@40055.4]
  assign _T_95111 = _T_94225 ? 16'h10 : _T_95110; // @[Mux.scala 31:69:@40056.4]
  assign _T_95112 = _T_94222 ? 16'h8 : _T_95111; // @[Mux.scala 31:69:@40057.4]
  assign _T_95113 = _T_94219 ? 16'h4 : _T_95112; // @[Mux.scala 31:69:@40058.4]
  assign _T_95114 = _T_94216 ? 16'h2 : _T_95113; // @[Mux.scala 31:69:@40059.4]
  assign _T_95115 = _T_94213 ? 16'h1 : _T_95114; // @[Mux.scala 31:69:@40060.4]
  assign _T_95116 = _T_95115[0]; // @[OneHot.scala 66:30:@40061.4]
  assign _T_95117 = _T_95115[1]; // @[OneHot.scala 66:30:@40062.4]
  assign _T_95118 = _T_95115[2]; // @[OneHot.scala 66:30:@40063.4]
  assign _T_95119 = _T_95115[3]; // @[OneHot.scala 66:30:@40064.4]
  assign _T_95120 = _T_95115[4]; // @[OneHot.scala 66:30:@40065.4]
  assign _T_95121 = _T_95115[5]; // @[OneHot.scala 66:30:@40066.4]
  assign _T_95122 = _T_95115[6]; // @[OneHot.scala 66:30:@40067.4]
  assign _T_95123 = _T_95115[7]; // @[OneHot.scala 66:30:@40068.4]
  assign _T_95124 = _T_95115[8]; // @[OneHot.scala 66:30:@40069.4]
  assign _T_95125 = _T_95115[9]; // @[OneHot.scala 66:30:@40070.4]
  assign _T_95126 = _T_95115[10]; // @[OneHot.scala 66:30:@40071.4]
  assign _T_95127 = _T_95115[11]; // @[OneHot.scala 66:30:@40072.4]
  assign _T_95128 = _T_95115[12]; // @[OneHot.scala 66:30:@40073.4]
  assign _T_95129 = _T_95115[13]; // @[OneHot.scala 66:30:@40074.4]
  assign _T_95130 = _T_95115[14]; // @[OneHot.scala 66:30:@40075.4]
  assign _T_95131 = _T_95115[15]; // @[OneHot.scala 66:30:@40076.4]
  assign _T_95172 = _T_94213 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40094.4]
  assign _T_95173 = _T_94210 ? 16'h4000 : _T_95172; // @[Mux.scala 31:69:@40095.4]
  assign _T_95174 = _T_94207 ? 16'h2000 : _T_95173; // @[Mux.scala 31:69:@40096.4]
  assign _T_95175 = _T_94204 ? 16'h1000 : _T_95174; // @[Mux.scala 31:69:@40097.4]
  assign _T_95176 = _T_94201 ? 16'h800 : _T_95175; // @[Mux.scala 31:69:@40098.4]
  assign _T_95177 = _T_94198 ? 16'h400 : _T_95176; // @[Mux.scala 31:69:@40099.4]
  assign _T_95178 = _T_94195 ? 16'h200 : _T_95177; // @[Mux.scala 31:69:@40100.4]
  assign _T_95179 = _T_94192 ? 16'h100 : _T_95178; // @[Mux.scala 31:69:@40101.4]
  assign _T_95180 = _T_94189 ? 16'h80 : _T_95179; // @[Mux.scala 31:69:@40102.4]
  assign _T_95181 = _T_94186 ? 16'h40 : _T_95180; // @[Mux.scala 31:69:@40103.4]
  assign _T_95182 = _T_94183 ? 16'h20 : _T_95181; // @[Mux.scala 31:69:@40104.4]
  assign _T_95183 = _T_94180 ? 16'h10 : _T_95182; // @[Mux.scala 31:69:@40105.4]
  assign _T_95184 = _T_94225 ? 16'h8 : _T_95183; // @[Mux.scala 31:69:@40106.4]
  assign _T_95185 = _T_94222 ? 16'h4 : _T_95184; // @[Mux.scala 31:69:@40107.4]
  assign _T_95186 = _T_94219 ? 16'h2 : _T_95185; // @[Mux.scala 31:69:@40108.4]
  assign _T_95187 = _T_94216 ? 16'h1 : _T_95186; // @[Mux.scala 31:69:@40109.4]
  assign _T_95188 = _T_95187[0]; // @[OneHot.scala 66:30:@40110.4]
  assign _T_95189 = _T_95187[1]; // @[OneHot.scala 66:30:@40111.4]
  assign _T_95190 = _T_95187[2]; // @[OneHot.scala 66:30:@40112.4]
  assign _T_95191 = _T_95187[3]; // @[OneHot.scala 66:30:@40113.4]
  assign _T_95192 = _T_95187[4]; // @[OneHot.scala 66:30:@40114.4]
  assign _T_95193 = _T_95187[5]; // @[OneHot.scala 66:30:@40115.4]
  assign _T_95194 = _T_95187[6]; // @[OneHot.scala 66:30:@40116.4]
  assign _T_95195 = _T_95187[7]; // @[OneHot.scala 66:30:@40117.4]
  assign _T_95196 = _T_95187[8]; // @[OneHot.scala 66:30:@40118.4]
  assign _T_95197 = _T_95187[9]; // @[OneHot.scala 66:30:@40119.4]
  assign _T_95198 = _T_95187[10]; // @[OneHot.scala 66:30:@40120.4]
  assign _T_95199 = _T_95187[11]; // @[OneHot.scala 66:30:@40121.4]
  assign _T_95200 = _T_95187[12]; // @[OneHot.scala 66:30:@40122.4]
  assign _T_95201 = _T_95187[13]; // @[OneHot.scala 66:30:@40123.4]
  assign _T_95202 = _T_95187[14]; // @[OneHot.scala 66:30:@40124.4]
  assign _T_95203 = _T_95187[15]; // @[OneHot.scala 66:30:@40125.4]
  assign _T_95244 = _T_94216 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40143.4]
  assign _T_95245 = _T_94213 ? 16'h4000 : _T_95244; // @[Mux.scala 31:69:@40144.4]
  assign _T_95246 = _T_94210 ? 16'h2000 : _T_95245; // @[Mux.scala 31:69:@40145.4]
  assign _T_95247 = _T_94207 ? 16'h1000 : _T_95246; // @[Mux.scala 31:69:@40146.4]
  assign _T_95248 = _T_94204 ? 16'h800 : _T_95247; // @[Mux.scala 31:69:@40147.4]
  assign _T_95249 = _T_94201 ? 16'h400 : _T_95248; // @[Mux.scala 31:69:@40148.4]
  assign _T_95250 = _T_94198 ? 16'h200 : _T_95249; // @[Mux.scala 31:69:@40149.4]
  assign _T_95251 = _T_94195 ? 16'h100 : _T_95250; // @[Mux.scala 31:69:@40150.4]
  assign _T_95252 = _T_94192 ? 16'h80 : _T_95251; // @[Mux.scala 31:69:@40151.4]
  assign _T_95253 = _T_94189 ? 16'h40 : _T_95252; // @[Mux.scala 31:69:@40152.4]
  assign _T_95254 = _T_94186 ? 16'h20 : _T_95253; // @[Mux.scala 31:69:@40153.4]
  assign _T_95255 = _T_94183 ? 16'h10 : _T_95254; // @[Mux.scala 31:69:@40154.4]
  assign _T_95256 = _T_94180 ? 16'h8 : _T_95255; // @[Mux.scala 31:69:@40155.4]
  assign _T_95257 = _T_94225 ? 16'h4 : _T_95256; // @[Mux.scala 31:69:@40156.4]
  assign _T_95258 = _T_94222 ? 16'h2 : _T_95257; // @[Mux.scala 31:69:@40157.4]
  assign _T_95259 = _T_94219 ? 16'h1 : _T_95258; // @[Mux.scala 31:69:@40158.4]
  assign _T_95260 = _T_95259[0]; // @[OneHot.scala 66:30:@40159.4]
  assign _T_95261 = _T_95259[1]; // @[OneHot.scala 66:30:@40160.4]
  assign _T_95262 = _T_95259[2]; // @[OneHot.scala 66:30:@40161.4]
  assign _T_95263 = _T_95259[3]; // @[OneHot.scala 66:30:@40162.4]
  assign _T_95264 = _T_95259[4]; // @[OneHot.scala 66:30:@40163.4]
  assign _T_95265 = _T_95259[5]; // @[OneHot.scala 66:30:@40164.4]
  assign _T_95266 = _T_95259[6]; // @[OneHot.scala 66:30:@40165.4]
  assign _T_95267 = _T_95259[7]; // @[OneHot.scala 66:30:@40166.4]
  assign _T_95268 = _T_95259[8]; // @[OneHot.scala 66:30:@40167.4]
  assign _T_95269 = _T_95259[9]; // @[OneHot.scala 66:30:@40168.4]
  assign _T_95270 = _T_95259[10]; // @[OneHot.scala 66:30:@40169.4]
  assign _T_95271 = _T_95259[11]; // @[OneHot.scala 66:30:@40170.4]
  assign _T_95272 = _T_95259[12]; // @[OneHot.scala 66:30:@40171.4]
  assign _T_95273 = _T_95259[13]; // @[OneHot.scala 66:30:@40172.4]
  assign _T_95274 = _T_95259[14]; // @[OneHot.scala 66:30:@40173.4]
  assign _T_95275 = _T_95259[15]; // @[OneHot.scala 66:30:@40174.4]
  assign _T_95316 = _T_94219 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40192.4]
  assign _T_95317 = _T_94216 ? 16'h4000 : _T_95316; // @[Mux.scala 31:69:@40193.4]
  assign _T_95318 = _T_94213 ? 16'h2000 : _T_95317; // @[Mux.scala 31:69:@40194.4]
  assign _T_95319 = _T_94210 ? 16'h1000 : _T_95318; // @[Mux.scala 31:69:@40195.4]
  assign _T_95320 = _T_94207 ? 16'h800 : _T_95319; // @[Mux.scala 31:69:@40196.4]
  assign _T_95321 = _T_94204 ? 16'h400 : _T_95320; // @[Mux.scala 31:69:@40197.4]
  assign _T_95322 = _T_94201 ? 16'h200 : _T_95321; // @[Mux.scala 31:69:@40198.4]
  assign _T_95323 = _T_94198 ? 16'h100 : _T_95322; // @[Mux.scala 31:69:@40199.4]
  assign _T_95324 = _T_94195 ? 16'h80 : _T_95323; // @[Mux.scala 31:69:@40200.4]
  assign _T_95325 = _T_94192 ? 16'h40 : _T_95324; // @[Mux.scala 31:69:@40201.4]
  assign _T_95326 = _T_94189 ? 16'h20 : _T_95325; // @[Mux.scala 31:69:@40202.4]
  assign _T_95327 = _T_94186 ? 16'h10 : _T_95326; // @[Mux.scala 31:69:@40203.4]
  assign _T_95328 = _T_94183 ? 16'h8 : _T_95327; // @[Mux.scala 31:69:@40204.4]
  assign _T_95329 = _T_94180 ? 16'h4 : _T_95328; // @[Mux.scala 31:69:@40205.4]
  assign _T_95330 = _T_94225 ? 16'h2 : _T_95329; // @[Mux.scala 31:69:@40206.4]
  assign _T_95331 = _T_94222 ? 16'h1 : _T_95330; // @[Mux.scala 31:69:@40207.4]
  assign _T_95332 = _T_95331[0]; // @[OneHot.scala 66:30:@40208.4]
  assign _T_95333 = _T_95331[1]; // @[OneHot.scala 66:30:@40209.4]
  assign _T_95334 = _T_95331[2]; // @[OneHot.scala 66:30:@40210.4]
  assign _T_95335 = _T_95331[3]; // @[OneHot.scala 66:30:@40211.4]
  assign _T_95336 = _T_95331[4]; // @[OneHot.scala 66:30:@40212.4]
  assign _T_95337 = _T_95331[5]; // @[OneHot.scala 66:30:@40213.4]
  assign _T_95338 = _T_95331[6]; // @[OneHot.scala 66:30:@40214.4]
  assign _T_95339 = _T_95331[7]; // @[OneHot.scala 66:30:@40215.4]
  assign _T_95340 = _T_95331[8]; // @[OneHot.scala 66:30:@40216.4]
  assign _T_95341 = _T_95331[9]; // @[OneHot.scala 66:30:@40217.4]
  assign _T_95342 = _T_95331[10]; // @[OneHot.scala 66:30:@40218.4]
  assign _T_95343 = _T_95331[11]; // @[OneHot.scala 66:30:@40219.4]
  assign _T_95344 = _T_95331[12]; // @[OneHot.scala 66:30:@40220.4]
  assign _T_95345 = _T_95331[13]; // @[OneHot.scala 66:30:@40221.4]
  assign _T_95346 = _T_95331[14]; // @[OneHot.scala 66:30:@40222.4]
  assign _T_95347 = _T_95331[15]; // @[OneHot.scala 66:30:@40223.4]
  assign _T_95388 = _T_94222 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40241.4]
  assign _T_95389 = _T_94219 ? 16'h4000 : _T_95388; // @[Mux.scala 31:69:@40242.4]
  assign _T_95390 = _T_94216 ? 16'h2000 : _T_95389; // @[Mux.scala 31:69:@40243.4]
  assign _T_95391 = _T_94213 ? 16'h1000 : _T_95390; // @[Mux.scala 31:69:@40244.4]
  assign _T_95392 = _T_94210 ? 16'h800 : _T_95391; // @[Mux.scala 31:69:@40245.4]
  assign _T_95393 = _T_94207 ? 16'h400 : _T_95392; // @[Mux.scala 31:69:@40246.4]
  assign _T_95394 = _T_94204 ? 16'h200 : _T_95393; // @[Mux.scala 31:69:@40247.4]
  assign _T_95395 = _T_94201 ? 16'h100 : _T_95394; // @[Mux.scala 31:69:@40248.4]
  assign _T_95396 = _T_94198 ? 16'h80 : _T_95395; // @[Mux.scala 31:69:@40249.4]
  assign _T_95397 = _T_94195 ? 16'h40 : _T_95396; // @[Mux.scala 31:69:@40250.4]
  assign _T_95398 = _T_94192 ? 16'h20 : _T_95397; // @[Mux.scala 31:69:@40251.4]
  assign _T_95399 = _T_94189 ? 16'h10 : _T_95398; // @[Mux.scala 31:69:@40252.4]
  assign _T_95400 = _T_94186 ? 16'h8 : _T_95399; // @[Mux.scala 31:69:@40253.4]
  assign _T_95401 = _T_94183 ? 16'h4 : _T_95400; // @[Mux.scala 31:69:@40254.4]
  assign _T_95402 = _T_94180 ? 16'h2 : _T_95401; // @[Mux.scala 31:69:@40255.4]
  assign _T_95403 = _T_94225 ? 16'h1 : _T_95402; // @[Mux.scala 31:69:@40256.4]
  assign _T_95404 = _T_95403[0]; // @[OneHot.scala 66:30:@40257.4]
  assign _T_95405 = _T_95403[1]; // @[OneHot.scala 66:30:@40258.4]
  assign _T_95406 = _T_95403[2]; // @[OneHot.scala 66:30:@40259.4]
  assign _T_95407 = _T_95403[3]; // @[OneHot.scala 66:30:@40260.4]
  assign _T_95408 = _T_95403[4]; // @[OneHot.scala 66:30:@40261.4]
  assign _T_95409 = _T_95403[5]; // @[OneHot.scala 66:30:@40262.4]
  assign _T_95410 = _T_95403[6]; // @[OneHot.scala 66:30:@40263.4]
  assign _T_95411 = _T_95403[7]; // @[OneHot.scala 66:30:@40264.4]
  assign _T_95412 = _T_95403[8]; // @[OneHot.scala 66:30:@40265.4]
  assign _T_95413 = _T_95403[9]; // @[OneHot.scala 66:30:@40266.4]
  assign _T_95414 = _T_95403[10]; // @[OneHot.scala 66:30:@40267.4]
  assign _T_95415 = _T_95403[11]; // @[OneHot.scala 66:30:@40268.4]
  assign _T_95416 = _T_95403[12]; // @[OneHot.scala 66:30:@40269.4]
  assign _T_95417 = _T_95403[13]; // @[OneHot.scala 66:30:@40270.4]
  assign _T_95418 = _T_95403[14]; // @[OneHot.scala 66:30:@40271.4]
  assign _T_95419 = _T_95403[15]; // @[OneHot.scala 66:30:@40272.4]
  assign _T_95484 = {_T_94331,_T_94330,_T_94329,_T_94328,_T_94327,_T_94326,_T_94325,_T_94324}; // @[Mux.scala 19:72:@40296.4]
  assign _T_95492 = {_T_94339,_T_94338,_T_94337,_T_94336,_T_94335,_T_94334,_T_94333,_T_94332,_T_95484}; // @[Mux.scala 19:72:@40304.4]
  assign _T_95494 = _T_90400 ? _T_95492 : 16'h0; // @[Mux.scala 19:72:@40305.4]
  assign _T_95501 = {_T_94402,_T_94401,_T_94400,_T_94399,_T_94398,_T_94397,_T_94396,_T_94411}; // @[Mux.scala 19:72:@40312.4]
  assign _T_95509 = {_T_94410,_T_94409,_T_94408,_T_94407,_T_94406,_T_94405,_T_94404,_T_94403,_T_95501}; // @[Mux.scala 19:72:@40320.4]
  assign _T_95511 = _T_90401 ? _T_95509 : 16'h0; // @[Mux.scala 19:72:@40321.4]
  assign _T_95518 = {_T_94473,_T_94472,_T_94471,_T_94470,_T_94469,_T_94468,_T_94483,_T_94482}; // @[Mux.scala 19:72:@40328.4]
  assign _T_95526 = {_T_94481,_T_94480,_T_94479,_T_94478,_T_94477,_T_94476,_T_94475,_T_94474,_T_95518}; // @[Mux.scala 19:72:@40336.4]
  assign _T_95528 = _T_90402 ? _T_95526 : 16'h0; // @[Mux.scala 19:72:@40337.4]
  assign _T_95535 = {_T_94544,_T_94543,_T_94542,_T_94541,_T_94540,_T_94555,_T_94554,_T_94553}; // @[Mux.scala 19:72:@40344.4]
  assign _T_95543 = {_T_94552,_T_94551,_T_94550,_T_94549,_T_94548,_T_94547,_T_94546,_T_94545,_T_95535}; // @[Mux.scala 19:72:@40352.4]
  assign _T_95545 = _T_90403 ? _T_95543 : 16'h0; // @[Mux.scala 19:72:@40353.4]
  assign _T_95552 = {_T_94615,_T_94614,_T_94613,_T_94612,_T_94627,_T_94626,_T_94625,_T_94624}; // @[Mux.scala 19:72:@40360.4]
  assign _T_95560 = {_T_94623,_T_94622,_T_94621,_T_94620,_T_94619,_T_94618,_T_94617,_T_94616,_T_95552}; // @[Mux.scala 19:72:@40368.4]
  assign _T_95562 = _T_90404 ? _T_95560 : 16'h0; // @[Mux.scala 19:72:@40369.4]
  assign _T_95569 = {_T_94686,_T_94685,_T_94684,_T_94699,_T_94698,_T_94697,_T_94696,_T_94695}; // @[Mux.scala 19:72:@40376.4]
  assign _T_95577 = {_T_94694,_T_94693,_T_94692,_T_94691,_T_94690,_T_94689,_T_94688,_T_94687,_T_95569}; // @[Mux.scala 19:72:@40384.4]
  assign _T_95579 = _T_90405 ? _T_95577 : 16'h0; // @[Mux.scala 19:72:@40385.4]
  assign _T_95586 = {_T_94757,_T_94756,_T_94771,_T_94770,_T_94769,_T_94768,_T_94767,_T_94766}; // @[Mux.scala 19:72:@40392.4]
  assign _T_95594 = {_T_94765,_T_94764,_T_94763,_T_94762,_T_94761,_T_94760,_T_94759,_T_94758,_T_95586}; // @[Mux.scala 19:72:@40400.4]
  assign _T_95596 = _T_90406 ? _T_95594 : 16'h0; // @[Mux.scala 19:72:@40401.4]
  assign _T_95603 = {_T_94828,_T_94843,_T_94842,_T_94841,_T_94840,_T_94839,_T_94838,_T_94837}; // @[Mux.scala 19:72:@40408.4]
  assign _T_95611 = {_T_94836,_T_94835,_T_94834,_T_94833,_T_94832,_T_94831,_T_94830,_T_94829,_T_95603}; // @[Mux.scala 19:72:@40416.4]
  assign _T_95613 = _T_90407 ? _T_95611 : 16'h0; // @[Mux.scala 19:72:@40417.4]
  assign _T_95620 = {_T_94915,_T_94914,_T_94913,_T_94912,_T_94911,_T_94910,_T_94909,_T_94908}; // @[Mux.scala 19:72:@40424.4]
  assign _T_95628 = {_T_94907,_T_94906,_T_94905,_T_94904,_T_94903,_T_94902,_T_94901,_T_94900,_T_95620}; // @[Mux.scala 19:72:@40432.4]
  assign _T_95630 = _T_90408 ? _T_95628 : 16'h0; // @[Mux.scala 19:72:@40433.4]
  assign _T_95637 = {_T_94986,_T_94985,_T_94984,_T_94983,_T_94982,_T_94981,_T_94980,_T_94979}; // @[Mux.scala 19:72:@40440.4]
  assign _T_95645 = {_T_94978,_T_94977,_T_94976,_T_94975,_T_94974,_T_94973,_T_94972,_T_94987,_T_95637}; // @[Mux.scala 19:72:@40448.4]
  assign _T_95647 = _T_90409 ? _T_95645 : 16'h0; // @[Mux.scala 19:72:@40449.4]
  assign _T_95654 = {_T_95057,_T_95056,_T_95055,_T_95054,_T_95053,_T_95052,_T_95051,_T_95050}; // @[Mux.scala 19:72:@40456.4]
  assign _T_95662 = {_T_95049,_T_95048,_T_95047,_T_95046,_T_95045,_T_95044,_T_95059,_T_95058,_T_95654}; // @[Mux.scala 19:72:@40464.4]
  assign _T_95664 = _T_90410 ? _T_95662 : 16'h0; // @[Mux.scala 19:72:@40465.4]
  assign _T_95671 = {_T_95128,_T_95127,_T_95126,_T_95125,_T_95124,_T_95123,_T_95122,_T_95121}; // @[Mux.scala 19:72:@40472.4]
  assign _T_95679 = {_T_95120,_T_95119,_T_95118,_T_95117,_T_95116,_T_95131,_T_95130,_T_95129,_T_95671}; // @[Mux.scala 19:72:@40480.4]
  assign _T_95681 = _T_90411 ? _T_95679 : 16'h0; // @[Mux.scala 19:72:@40481.4]
  assign _T_95688 = {_T_95199,_T_95198,_T_95197,_T_95196,_T_95195,_T_95194,_T_95193,_T_95192}; // @[Mux.scala 19:72:@40488.4]
  assign _T_95696 = {_T_95191,_T_95190,_T_95189,_T_95188,_T_95203,_T_95202,_T_95201,_T_95200,_T_95688}; // @[Mux.scala 19:72:@40496.4]
  assign _T_95698 = _T_90412 ? _T_95696 : 16'h0; // @[Mux.scala 19:72:@40497.4]
  assign _T_95705 = {_T_95270,_T_95269,_T_95268,_T_95267,_T_95266,_T_95265,_T_95264,_T_95263}; // @[Mux.scala 19:72:@40504.4]
  assign _T_95713 = {_T_95262,_T_95261,_T_95260,_T_95275,_T_95274,_T_95273,_T_95272,_T_95271,_T_95705}; // @[Mux.scala 19:72:@40512.4]
  assign _T_95715 = _T_90413 ? _T_95713 : 16'h0; // @[Mux.scala 19:72:@40513.4]
  assign _T_95722 = {_T_95341,_T_95340,_T_95339,_T_95338,_T_95337,_T_95336,_T_95335,_T_95334}; // @[Mux.scala 19:72:@40520.4]
  assign _T_95730 = {_T_95333,_T_95332,_T_95347,_T_95346,_T_95345,_T_95344,_T_95343,_T_95342,_T_95722}; // @[Mux.scala 19:72:@40528.4]
  assign _T_95732 = _T_90414 ? _T_95730 : 16'h0; // @[Mux.scala 19:72:@40529.4]
  assign _T_95739 = {_T_95412,_T_95411,_T_95410,_T_95409,_T_95408,_T_95407,_T_95406,_T_95405}; // @[Mux.scala 19:72:@40536.4]
  assign _T_95747 = {_T_95404,_T_95419,_T_95418,_T_95417,_T_95416,_T_95415,_T_95414,_T_95413,_T_95739}; // @[Mux.scala 19:72:@40544.4]
  assign _T_95749 = _T_90415 ? _T_95747 : 16'h0; // @[Mux.scala 19:72:@40545.4]
  assign _T_95750 = _T_95494 | _T_95511; // @[Mux.scala 19:72:@40546.4]
  assign _T_95751 = _T_95750 | _T_95528; // @[Mux.scala 19:72:@40547.4]
  assign _T_95752 = _T_95751 | _T_95545; // @[Mux.scala 19:72:@40548.4]
  assign _T_95753 = _T_95752 | _T_95562; // @[Mux.scala 19:72:@40549.4]
  assign _T_95754 = _T_95753 | _T_95579; // @[Mux.scala 19:72:@40550.4]
  assign _T_95755 = _T_95754 | _T_95596; // @[Mux.scala 19:72:@40551.4]
  assign _T_95756 = _T_95755 | _T_95613; // @[Mux.scala 19:72:@40552.4]
  assign _T_95757 = _T_95756 | _T_95630; // @[Mux.scala 19:72:@40553.4]
  assign _T_95758 = _T_95757 | _T_95647; // @[Mux.scala 19:72:@40554.4]
  assign _T_95759 = _T_95758 | _T_95664; // @[Mux.scala 19:72:@40555.4]
  assign _T_95760 = _T_95759 | _T_95681; // @[Mux.scala 19:72:@40556.4]
  assign _T_95761 = _T_95760 | _T_95698; // @[Mux.scala 19:72:@40557.4]
  assign _T_95762 = _T_95761 | _T_95715; // @[Mux.scala 19:72:@40558.4]
  assign _T_95763 = _T_95762 | _T_95732; // @[Mux.scala 19:72:@40559.4]
  assign _T_95764 = _T_95763 | _T_95749; // @[Mux.scala 19:72:@40560.4]
  assign inputPriorityPorts_0_0 = _T_95764[0]; // @[Mux.scala 19:72:@40564.4]
  assign inputPriorityPorts_0_1 = _T_95764[1]; // @[Mux.scala 19:72:@40566.4]
  assign inputPriorityPorts_0_2 = _T_95764[2]; // @[Mux.scala 19:72:@40568.4]
  assign inputPriorityPorts_0_3 = _T_95764[3]; // @[Mux.scala 19:72:@40570.4]
  assign inputPriorityPorts_0_4 = _T_95764[4]; // @[Mux.scala 19:72:@40572.4]
  assign inputPriorityPorts_0_5 = _T_95764[5]; // @[Mux.scala 19:72:@40574.4]
  assign inputPriorityPorts_0_6 = _T_95764[6]; // @[Mux.scala 19:72:@40576.4]
  assign inputPriorityPorts_0_7 = _T_95764[7]; // @[Mux.scala 19:72:@40578.4]
  assign inputPriorityPorts_0_8 = _T_95764[8]; // @[Mux.scala 19:72:@40580.4]
  assign inputPriorityPorts_0_9 = _T_95764[9]; // @[Mux.scala 19:72:@40582.4]
  assign inputPriorityPorts_0_10 = _T_95764[10]; // @[Mux.scala 19:72:@40584.4]
  assign inputPriorityPorts_0_11 = _T_95764[11]; // @[Mux.scala 19:72:@40586.4]
  assign inputPriorityPorts_0_12 = _T_95764[12]; // @[Mux.scala 19:72:@40588.4]
  assign inputPriorityPorts_0_13 = _T_95764[13]; // @[Mux.scala 19:72:@40590.4]
  assign inputPriorityPorts_0_14 = _T_95764[14]; // @[Mux.scala 19:72:@40592.4]
  assign inputPriorityPorts_0_15 = _T_95764[15]; // @[Mux.scala 19:72:@40594.4]
  assign _T_95966 = entriesPorts_0_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40648.4]
  assign _T_95967 = entriesPorts_0_14 ? 16'h4000 : _T_95966; // @[Mux.scala 31:69:@40649.4]
  assign _T_95968 = entriesPorts_0_13 ? 16'h2000 : _T_95967; // @[Mux.scala 31:69:@40650.4]
  assign _T_95969 = entriesPorts_0_12 ? 16'h1000 : _T_95968; // @[Mux.scala 31:69:@40651.4]
  assign _T_95970 = entriesPorts_0_11 ? 16'h800 : _T_95969; // @[Mux.scala 31:69:@40652.4]
  assign _T_95971 = entriesPorts_0_10 ? 16'h400 : _T_95970; // @[Mux.scala 31:69:@40653.4]
  assign _T_95972 = entriesPorts_0_9 ? 16'h200 : _T_95971; // @[Mux.scala 31:69:@40654.4]
  assign _T_95973 = entriesPorts_0_8 ? 16'h100 : _T_95972; // @[Mux.scala 31:69:@40655.4]
  assign _T_95974 = entriesPorts_0_7 ? 16'h80 : _T_95973; // @[Mux.scala 31:69:@40656.4]
  assign _T_95975 = entriesPorts_0_6 ? 16'h40 : _T_95974; // @[Mux.scala 31:69:@40657.4]
  assign _T_95976 = entriesPorts_0_5 ? 16'h20 : _T_95975; // @[Mux.scala 31:69:@40658.4]
  assign _T_95977 = entriesPorts_0_4 ? 16'h10 : _T_95976; // @[Mux.scala 31:69:@40659.4]
  assign _T_95978 = entriesPorts_0_3 ? 16'h8 : _T_95977; // @[Mux.scala 31:69:@40660.4]
  assign _T_95979 = entriesPorts_0_2 ? 16'h4 : _T_95978; // @[Mux.scala 31:69:@40661.4]
  assign _T_95980 = entriesPorts_0_1 ? 16'h2 : _T_95979; // @[Mux.scala 31:69:@40662.4]
  assign _T_95981 = entriesPorts_0_0 ? 16'h1 : _T_95980; // @[Mux.scala 31:69:@40663.4]
  assign _T_95982 = _T_95981[0]; // @[OneHot.scala 66:30:@40664.4]
  assign _T_95983 = _T_95981[1]; // @[OneHot.scala 66:30:@40665.4]
  assign _T_95984 = _T_95981[2]; // @[OneHot.scala 66:30:@40666.4]
  assign _T_95985 = _T_95981[3]; // @[OneHot.scala 66:30:@40667.4]
  assign _T_95986 = _T_95981[4]; // @[OneHot.scala 66:30:@40668.4]
  assign _T_95987 = _T_95981[5]; // @[OneHot.scala 66:30:@40669.4]
  assign _T_95988 = _T_95981[6]; // @[OneHot.scala 66:30:@40670.4]
  assign _T_95989 = _T_95981[7]; // @[OneHot.scala 66:30:@40671.4]
  assign _T_95990 = _T_95981[8]; // @[OneHot.scala 66:30:@40672.4]
  assign _T_95991 = _T_95981[9]; // @[OneHot.scala 66:30:@40673.4]
  assign _T_95992 = _T_95981[10]; // @[OneHot.scala 66:30:@40674.4]
  assign _T_95993 = _T_95981[11]; // @[OneHot.scala 66:30:@40675.4]
  assign _T_95994 = _T_95981[12]; // @[OneHot.scala 66:30:@40676.4]
  assign _T_95995 = _T_95981[13]; // @[OneHot.scala 66:30:@40677.4]
  assign _T_95996 = _T_95981[14]; // @[OneHot.scala 66:30:@40678.4]
  assign _T_95997 = _T_95981[15]; // @[OneHot.scala 66:30:@40679.4]
  assign _T_96038 = entriesPorts_0_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40697.4]
  assign _T_96039 = entriesPorts_0_15 ? 16'h4000 : _T_96038; // @[Mux.scala 31:69:@40698.4]
  assign _T_96040 = entriesPorts_0_14 ? 16'h2000 : _T_96039; // @[Mux.scala 31:69:@40699.4]
  assign _T_96041 = entriesPorts_0_13 ? 16'h1000 : _T_96040; // @[Mux.scala 31:69:@40700.4]
  assign _T_96042 = entriesPorts_0_12 ? 16'h800 : _T_96041; // @[Mux.scala 31:69:@40701.4]
  assign _T_96043 = entriesPorts_0_11 ? 16'h400 : _T_96042; // @[Mux.scala 31:69:@40702.4]
  assign _T_96044 = entriesPorts_0_10 ? 16'h200 : _T_96043; // @[Mux.scala 31:69:@40703.4]
  assign _T_96045 = entriesPorts_0_9 ? 16'h100 : _T_96044; // @[Mux.scala 31:69:@40704.4]
  assign _T_96046 = entriesPorts_0_8 ? 16'h80 : _T_96045; // @[Mux.scala 31:69:@40705.4]
  assign _T_96047 = entriesPorts_0_7 ? 16'h40 : _T_96046; // @[Mux.scala 31:69:@40706.4]
  assign _T_96048 = entriesPorts_0_6 ? 16'h20 : _T_96047; // @[Mux.scala 31:69:@40707.4]
  assign _T_96049 = entriesPorts_0_5 ? 16'h10 : _T_96048; // @[Mux.scala 31:69:@40708.4]
  assign _T_96050 = entriesPorts_0_4 ? 16'h8 : _T_96049; // @[Mux.scala 31:69:@40709.4]
  assign _T_96051 = entriesPorts_0_3 ? 16'h4 : _T_96050; // @[Mux.scala 31:69:@40710.4]
  assign _T_96052 = entriesPorts_0_2 ? 16'h2 : _T_96051; // @[Mux.scala 31:69:@40711.4]
  assign _T_96053 = entriesPorts_0_1 ? 16'h1 : _T_96052; // @[Mux.scala 31:69:@40712.4]
  assign _T_96054 = _T_96053[0]; // @[OneHot.scala 66:30:@40713.4]
  assign _T_96055 = _T_96053[1]; // @[OneHot.scala 66:30:@40714.4]
  assign _T_96056 = _T_96053[2]; // @[OneHot.scala 66:30:@40715.4]
  assign _T_96057 = _T_96053[3]; // @[OneHot.scala 66:30:@40716.4]
  assign _T_96058 = _T_96053[4]; // @[OneHot.scala 66:30:@40717.4]
  assign _T_96059 = _T_96053[5]; // @[OneHot.scala 66:30:@40718.4]
  assign _T_96060 = _T_96053[6]; // @[OneHot.scala 66:30:@40719.4]
  assign _T_96061 = _T_96053[7]; // @[OneHot.scala 66:30:@40720.4]
  assign _T_96062 = _T_96053[8]; // @[OneHot.scala 66:30:@40721.4]
  assign _T_96063 = _T_96053[9]; // @[OneHot.scala 66:30:@40722.4]
  assign _T_96064 = _T_96053[10]; // @[OneHot.scala 66:30:@40723.4]
  assign _T_96065 = _T_96053[11]; // @[OneHot.scala 66:30:@40724.4]
  assign _T_96066 = _T_96053[12]; // @[OneHot.scala 66:30:@40725.4]
  assign _T_96067 = _T_96053[13]; // @[OneHot.scala 66:30:@40726.4]
  assign _T_96068 = _T_96053[14]; // @[OneHot.scala 66:30:@40727.4]
  assign _T_96069 = _T_96053[15]; // @[OneHot.scala 66:30:@40728.4]
  assign _T_96110 = entriesPorts_0_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40746.4]
  assign _T_96111 = entriesPorts_0_0 ? 16'h4000 : _T_96110; // @[Mux.scala 31:69:@40747.4]
  assign _T_96112 = entriesPorts_0_15 ? 16'h2000 : _T_96111; // @[Mux.scala 31:69:@40748.4]
  assign _T_96113 = entriesPorts_0_14 ? 16'h1000 : _T_96112; // @[Mux.scala 31:69:@40749.4]
  assign _T_96114 = entriesPorts_0_13 ? 16'h800 : _T_96113; // @[Mux.scala 31:69:@40750.4]
  assign _T_96115 = entriesPorts_0_12 ? 16'h400 : _T_96114; // @[Mux.scala 31:69:@40751.4]
  assign _T_96116 = entriesPorts_0_11 ? 16'h200 : _T_96115; // @[Mux.scala 31:69:@40752.4]
  assign _T_96117 = entriesPorts_0_10 ? 16'h100 : _T_96116; // @[Mux.scala 31:69:@40753.4]
  assign _T_96118 = entriesPorts_0_9 ? 16'h80 : _T_96117; // @[Mux.scala 31:69:@40754.4]
  assign _T_96119 = entriesPorts_0_8 ? 16'h40 : _T_96118; // @[Mux.scala 31:69:@40755.4]
  assign _T_96120 = entriesPorts_0_7 ? 16'h20 : _T_96119; // @[Mux.scala 31:69:@40756.4]
  assign _T_96121 = entriesPorts_0_6 ? 16'h10 : _T_96120; // @[Mux.scala 31:69:@40757.4]
  assign _T_96122 = entriesPorts_0_5 ? 16'h8 : _T_96121; // @[Mux.scala 31:69:@40758.4]
  assign _T_96123 = entriesPorts_0_4 ? 16'h4 : _T_96122; // @[Mux.scala 31:69:@40759.4]
  assign _T_96124 = entriesPorts_0_3 ? 16'h2 : _T_96123; // @[Mux.scala 31:69:@40760.4]
  assign _T_96125 = entriesPorts_0_2 ? 16'h1 : _T_96124; // @[Mux.scala 31:69:@40761.4]
  assign _T_96126 = _T_96125[0]; // @[OneHot.scala 66:30:@40762.4]
  assign _T_96127 = _T_96125[1]; // @[OneHot.scala 66:30:@40763.4]
  assign _T_96128 = _T_96125[2]; // @[OneHot.scala 66:30:@40764.4]
  assign _T_96129 = _T_96125[3]; // @[OneHot.scala 66:30:@40765.4]
  assign _T_96130 = _T_96125[4]; // @[OneHot.scala 66:30:@40766.4]
  assign _T_96131 = _T_96125[5]; // @[OneHot.scala 66:30:@40767.4]
  assign _T_96132 = _T_96125[6]; // @[OneHot.scala 66:30:@40768.4]
  assign _T_96133 = _T_96125[7]; // @[OneHot.scala 66:30:@40769.4]
  assign _T_96134 = _T_96125[8]; // @[OneHot.scala 66:30:@40770.4]
  assign _T_96135 = _T_96125[9]; // @[OneHot.scala 66:30:@40771.4]
  assign _T_96136 = _T_96125[10]; // @[OneHot.scala 66:30:@40772.4]
  assign _T_96137 = _T_96125[11]; // @[OneHot.scala 66:30:@40773.4]
  assign _T_96138 = _T_96125[12]; // @[OneHot.scala 66:30:@40774.4]
  assign _T_96139 = _T_96125[13]; // @[OneHot.scala 66:30:@40775.4]
  assign _T_96140 = _T_96125[14]; // @[OneHot.scala 66:30:@40776.4]
  assign _T_96141 = _T_96125[15]; // @[OneHot.scala 66:30:@40777.4]
  assign _T_96182 = entriesPorts_0_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40795.4]
  assign _T_96183 = entriesPorts_0_1 ? 16'h4000 : _T_96182; // @[Mux.scala 31:69:@40796.4]
  assign _T_96184 = entriesPorts_0_0 ? 16'h2000 : _T_96183; // @[Mux.scala 31:69:@40797.4]
  assign _T_96185 = entriesPorts_0_15 ? 16'h1000 : _T_96184; // @[Mux.scala 31:69:@40798.4]
  assign _T_96186 = entriesPorts_0_14 ? 16'h800 : _T_96185; // @[Mux.scala 31:69:@40799.4]
  assign _T_96187 = entriesPorts_0_13 ? 16'h400 : _T_96186; // @[Mux.scala 31:69:@40800.4]
  assign _T_96188 = entriesPorts_0_12 ? 16'h200 : _T_96187; // @[Mux.scala 31:69:@40801.4]
  assign _T_96189 = entriesPorts_0_11 ? 16'h100 : _T_96188; // @[Mux.scala 31:69:@40802.4]
  assign _T_96190 = entriesPorts_0_10 ? 16'h80 : _T_96189; // @[Mux.scala 31:69:@40803.4]
  assign _T_96191 = entriesPorts_0_9 ? 16'h40 : _T_96190; // @[Mux.scala 31:69:@40804.4]
  assign _T_96192 = entriesPorts_0_8 ? 16'h20 : _T_96191; // @[Mux.scala 31:69:@40805.4]
  assign _T_96193 = entriesPorts_0_7 ? 16'h10 : _T_96192; // @[Mux.scala 31:69:@40806.4]
  assign _T_96194 = entriesPorts_0_6 ? 16'h8 : _T_96193; // @[Mux.scala 31:69:@40807.4]
  assign _T_96195 = entriesPorts_0_5 ? 16'h4 : _T_96194; // @[Mux.scala 31:69:@40808.4]
  assign _T_96196 = entriesPorts_0_4 ? 16'h2 : _T_96195; // @[Mux.scala 31:69:@40809.4]
  assign _T_96197 = entriesPorts_0_3 ? 16'h1 : _T_96196; // @[Mux.scala 31:69:@40810.4]
  assign _T_96198 = _T_96197[0]; // @[OneHot.scala 66:30:@40811.4]
  assign _T_96199 = _T_96197[1]; // @[OneHot.scala 66:30:@40812.4]
  assign _T_96200 = _T_96197[2]; // @[OneHot.scala 66:30:@40813.4]
  assign _T_96201 = _T_96197[3]; // @[OneHot.scala 66:30:@40814.4]
  assign _T_96202 = _T_96197[4]; // @[OneHot.scala 66:30:@40815.4]
  assign _T_96203 = _T_96197[5]; // @[OneHot.scala 66:30:@40816.4]
  assign _T_96204 = _T_96197[6]; // @[OneHot.scala 66:30:@40817.4]
  assign _T_96205 = _T_96197[7]; // @[OneHot.scala 66:30:@40818.4]
  assign _T_96206 = _T_96197[8]; // @[OneHot.scala 66:30:@40819.4]
  assign _T_96207 = _T_96197[9]; // @[OneHot.scala 66:30:@40820.4]
  assign _T_96208 = _T_96197[10]; // @[OneHot.scala 66:30:@40821.4]
  assign _T_96209 = _T_96197[11]; // @[OneHot.scala 66:30:@40822.4]
  assign _T_96210 = _T_96197[12]; // @[OneHot.scala 66:30:@40823.4]
  assign _T_96211 = _T_96197[13]; // @[OneHot.scala 66:30:@40824.4]
  assign _T_96212 = _T_96197[14]; // @[OneHot.scala 66:30:@40825.4]
  assign _T_96213 = _T_96197[15]; // @[OneHot.scala 66:30:@40826.4]
  assign _T_96254 = entriesPorts_0_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40844.4]
  assign _T_96255 = entriesPorts_0_2 ? 16'h4000 : _T_96254; // @[Mux.scala 31:69:@40845.4]
  assign _T_96256 = entriesPorts_0_1 ? 16'h2000 : _T_96255; // @[Mux.scala 31:69:@40846.4]
  assign _T_96257 = entriesPorts_0_0 ? 16'h1000 : _T_96256; // @[Mux.scala 31:69:@40847.4]
  assign _T_96258 = entriesPorts_0_15 ? 16'h800 : _T_96257; // @[Mux.scala 31:69:@40848.4]
  assign _T_96259 = entriesPorts_0_14 ? 16'h400 : _T_96258; // @[Mux.scala 31:69:@40849.4]
  assign _T_96260 = entriesPorts_0_13 ? 16'h200 : _T_96259; // @[Mux.scala 31:69:@40850.4]
  assign _T_96261 = entriesPorts_0_12 ? 16'h100 : _T_96260; // @[Mux.scala 31:69:@40851.4]
  assign _T_96262 = entriesPorts_0_11 ? 16'h80 : _T_96261; // @[Mux.scala 31:69:@40852.4]
  assign _T_96263 = entriesPorts_0_10 ? 16'h40 : _T_96262; // @[Mux.scala 31:69:@40853.4]
  assign _T_96264 = entriesPorts_0_9 ? 16'h20 : _T_96263; // @[Mux.scala 31:69:@40854.4]
  assign _T_96265 = entriesPorts_0_8 ? 16'h10 : _T_96264; // @[Mux.scala 31:69:@40855.4]
  assign _T_96266 = entriesPorts_0_7 ? 16'h8 : _T_96265; // @[Mux.scala 31:69:@40856.4]
  assign _T_96267 = entriesPorts_0_6 ? 16'h4 : _T_96266; // @[Mux.scala 31:69:@40857.4]
  assign _T_96268 = entriesPorts_0_5 ? 16'h2 : _T_96267; // @[Mux.scala 31:69:@40858.4]
  assign _T_96269 = entriesPorts_0_4 ? 16'h1 : _T_96268; // @[Mux.scala 31:69:@40859.4]
  assign _T_96270 = _T_96269[0]; // @[OneHot.scala 66:30:@40860.4]
  assign _T_96271 = _T_96269[1]; // @[OneHot.scala 66:30:@40861.4]
  assign _T_96272 = _T_96269[2]; // @[OneHot.scala 66:30:@40862.4]
  assign _T_96273 = _T_96269[3]; // @[OneHot.scala 66:30:@40863.4]
  assign _T_96274 = _T_96269[4]; // @[OneHot.scala 66:30:@40864.4]
  assign _T_96275 = _T_96269[5]; // @[OneHot.scala 66:30:@40865.4]
  assign _T_96276 = _T_96269[6]; // @[OneHot.scala 66:30:@40866.4]
  assign _T_96277 = _T_96269[7]; // @[OneHot.scala 66:30:@40867.4]
  assign _T_96278 = _T_96269[8]; // @[OneHot.scala 66:30:@40868.4]
  assign _T_96279 = _T_96269[9]; // @[OneHot.scala 66:30:@40869.4]
  assign _T_96280 = _T_96269[10]; // @[OneHot.scala 66:30:@40870.4]
  assign _T_96281 = _T_96269[11]; // @[OneHot.scala 66:30:@40871.4]
  assign _T_96282 = _T_96269[12]; // @[OneHot.scala 66:30:@40872.4]
  assign _T_96283 = _T_96269[13]; // @[OneHot.scala 66:30:@40873.4]
  assign _T_96284 = _T_96269[14]; // @[OneHot.scala 66:30:@40874.4]
  assign _T_96285 = _T_96269[15]; // @[OneHot.scala 66:30:@40875.4]
  assign _T_96326 = entriesPorts_0_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40893.4]
  assign _T_96327 = entriesPorts_0_3 ? 16'h4000 : _T_96326; // @[Mux.scala 31:69:@40894.4]
  assign _T_96328 = entriesPorts_0_2 ? 16'h2000 : _T_96327; // @[Mux.scala 31:69:@40895.4]
  assign _T_96329 = entriesPorts_0_1 ? 16'h1000 : _T_96328; // @[Mux.scala 31:69:@40896.4]
  assign _T_96330 = entriesPorts_0_0 ? 16'h800 : _T_96329; // @[Mux.scala 31:69:@40897.4]
  assign _T_96331 = entriesPorts_0_15 ? 16'h400 : _T_96330; // @[Mux.scala 31:69:@40898.4]
  assign _T_96332 = entriesPorts_0_14 ? 16'h200 : _T_96331; // @[Mux.scala 31:69:@40899.4]
  assign _T_96333 = entriesPorts_0_13 ? 16'h100 : _T_96332; // @[Mux.scala 31:69:@40900.4]
  assign _T_96334 = entriesPorts_0_12 ? 16'h80 : _T_96333; // @[Mux.scala 31:69:@40901.4]
  assign _T_96335 = entriesPorts_0_11 ? 16'h40 : _T_96334; // @[Mux.scala 31:69:@40902.4]
  assign _T_96336 = entriesPorts_0_10 ? 16'h20 : _T_96335; // @[Mux.scala 31:69:@40903.4]
  assign _T_96337 = entriesPorts_0_9 ? 16'h10 : _T_96336; // @[Mux.scala 31:69:@40904.4]
  assign _T_96338 = entriesPorts_0_8 ? 16'h8 : _T_96337; // @[Mux.scala 31:69:@40905.4]
  assign _T_96339 = entriesPorts_0_7 ? 16'h4 : _T_96338; // @[Mux.scala 31:69:@40906.4]
  assign _T_96340 = entriesPorts_0_6 ? 16'h2 : _T_96339; // @[Mux.scala 31:69:@40907.4]
  assign _T_96341 = entriesPorts_0_5 ? 16'h1 : _T_96340; // @[Mux.scala 31:69:@40908.4]
  assign _T_96342 = _T_96341[0]; // @[OneHot.scala 66:30:@40909.4]
  assign _T_96343 = _T_96341[1]; // @[OneHot.scala 66:30:@40910.4]
  assign _T_96344 = _T_96341[2]; // @[OneHot.scala 66:30:@40911.4]
  assign _T_96345 = _T_96341[3]; // @[OneHot.scala 66:30:@40912.4]
  assign _T_96346 = _T_96341[4]; // @[OneHot.scala 66:30:@40913.4]
  assign _T_96347 = _T_96341[5]; // @[OneHot.scala 66:30:@40914.4]
  assign _T_96348 = _T_96341[6]; // @[OneHot.scala 66:30:@40915.4]
  assign _T_96349 = _T_96341[7]; // @[OneHot.scala 66:30:@40916.4]
  assign _T_96350 = _T_96341[8]; // @[OneHot.scala 66:30:@40917.4]
  assign _T_96351 = _T_96341[9]; // @[OneHot.scala 66:30:@40918.4]
  assign _T_96352 = _T_96341[10]; // @[OneHot.scala 66:30:@40919.4]
  assign _T_96353 = _T_96341[11]; // @[OneHot.scala 66:30:@40920.4]
  assign _T_96354 = _T_96341[12]; // @[OneHot.scala 66:30:@40921.4]
  assign _T_96355 = _T_96341[13]; // @[OneHot.scala 66:30:@40922.4]
  assign _T_96356 = _T_96341[14]; // @[OneHot.scala 66:30:@40923.4]
  assign _T_96357 = _T_96341[15]; // @[OneHot.scala 66:30:@40924.4]
  assign _T_96398 = entriesPorts_0_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40942.4]
  assign _T_96399 = entriesPorts_0_4 ? 16'h4000 : _T_96398; // @[Mux.scala 31:69:@40943.4]
  assign _T_96400 = entriesPorts_0_3 ? 16'h2000 : _T_96399; // @[Mux.scala 31:69:@40944.4]
  assign _T_96401 = entriesPorts_0_2 ? 16'h1000 : _T_96400; // @[Mux.scala 31:69:@40945.4]
  assign _T_96402 = entriesPorts_0_1 ? 16'h800 : _T_96401; // @[Mux.scala 31:69:@40946.4]
  assign _T_96403 = entriesPorts_0_0 ? 16'h400 : _T_96402; // @[Mux.scala 31:69:@40947.4]
  assign _T_96404 = entriesPorts_0_15 ? 16'h200 : _T_96403; // @[Mux.scala 31:69:@40948.4]
  assign _T_96405 = entriesPorts_0_14 ? 16'h100 : _T_96404; // @[Mux.scala 31:69:@40949.4]
  assign _T_96406 = entriesPorts_0_13 ? 16'h80 : _T_96405; // @[Mux.scala 31:69:@40950.4]
  assign _T_96407 = entriesPorts_0_12 ? 16'h40 : _T_96406; // @[Mux.scala 31:69:@40951.4]
  assign _T_96408 = entriesPorts_0_11 ? 16'h20 : _T_96407; // @[Mux.scala 31:69:@40952.4]
  assign _T_96409 = entriesPorts_0_10 ? 16'h10 : _T_96408; // @[Mux.scala 31:69:@40953.4]
  assign _T_96410 = entriesPorts_0_9 ? 16'h8 : _T_96409; // @[Mux.scala 31:69:@40954.4]
  assign _T_96411 = entriesPorts_0_8 ? 16'h4 : _T_96410; // @[Mux.scala 31:69:@40955.4]
  assign _T_96412 = entriesPorts_0_7 ? 16'h2 : _T_96411; // @[Mux.scala 31:69:@40956.4]
  assign _T_96413 = entriesPorts_0_6 ? 16'h1 : _T_96412; // @[Mux.scala 31:69:@40957.4]
  assign _T_96414 = _T_96413[0]; // @[OneHot.scala 66:30:@40958.4]
  assign _T_96415 = _T_96413[1]; // @[OneHot.scala 66:30:@40959.4]
  assign _T_96416 = _T_96413[2]; // @[OneHot.scala 66:30:@40960.4]
  assign _T_96417 = _T_96413[3]; // @[OneHot.scala 66:30:@40961.4]
  assign _T_96418 = _T_96413[4]; // @[OneHot.scala 66:30:@40962.4]
  assign _T_96419 = _T_96413[5]; // @[OneHot.scala 66:30:@40963.4]
  assign _T_96420 = _T_96413[6]; // @[OneHot.scala 66:30:@40964.4]
  assign _T_96421 = _T_96413[7]; // @[OneHot.scala 66:30:@40965.4]
  assign _T_96422 = _T_96413[8]; // @[OneHot.scala 66:30:@40966.4]
  assign _T_96423 = _T_96413[9]; // @[OneHot.scala 66:30:@40967.4]
  assign _T_96424 = _T_96413[10]; // @[OneHot.scala 66:30:@40968.4]
  assign _T_96425 = _T_96413[11]; // @[OneHot.scala 66:30:@40969.4]
  assign _T_96426 = _T_96413[12]; // @[OneHot.scala 66:30:@40970.4]
  assign _T_96427 = _T_96413[13]; // @[OneHot.scala 66:30:@40971.4]
  assign _T_96428 = _T_96413[14]; // @[OneHot.scala 66:30:@40972.4]
  assign _T_96429 = _T_96413[15]; // @[OneHot.scala 66:30:@40973.4]
  assign _T_96470 = entriesPorts_0_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40991.4]
  assign _T_96471 = entriesPorts_0_5 ? 16'h4000 : _T_96470; // @[Mux.scala 31:69:@40992.4]
  assign _T_96472 = entriesPorts_0_4 ? 16'h2000 : _T_96471; // @[Mux.scala 31:69:@40993.4]
  assign _T_96473 = entriesPorts_0_3 ? 16'h1000 : _T_96472; // @[Mux.scala 31:69:@40994.4]
  assign _T_96474 = entriesPorts_0_2 ? 16'h800 : _T_96473; // @[Mux.scala 31:69:@40995.4]
  assign _T_96475 = entriesPorts_0_1 ? 16'h400 : _T_96474; // @[Mux.scala 31:69:@40996.4]
  assign _T_96476 = entriesPorts_0_0 ? 16'h200 : _T_96475; // @[Mux.scala 31:69:@40997.4]
  assign _T_96477 = entriesPorts_0_15 ? 16'h100 : _T_96476; // @[Mux.scala 31:69:@40998.4]
  assign _T_96478 = entriesPorts_0_14 ? 16'h80 : _T_96477; // @[Mux.scala 31:69:@40999.4]
  assign _T_96479 = entriesPorts_0_13 ? 16'h40 : _T_96478; // @[Mux.scala 31:69:@41000.4]
  assign _T_96480 = entriesPorts_0_12 ? 16'h20 : _T_96479; // @[Mux.scala 31:69:@41001.4]
  assign _T_96481 = entriesPorts_0_11 ? 16'h10 : _T_96480; // @[Mux.scala 31:69:@41002.4]
  assign _T_96482 = entriesPorts_0_10 ? 16'h8 : _T_96481; // @[Mux.scala 31:69:@41003.4]
  assign _T_96483 = entriesPorts_0_9 ? 16'h4 : _T_96482; // @[Mux.scala 31:69:@41004.4]
  assign _T_96484 = entriesPorts_0_8 ? 16'h2 : _T_96483; // @[Mux.scala 31:69:@41005.4]
  assign _T_96485 = entriesPorts_0_7 ? 16'h1 : _T_96484; // @[Mux.scala 31:69:@41006.4]
  assign _T_96486 = _T_96485[0]; // @[OneHot.scala 66:30:@41007.4]
  assign _T_96487 = _T_96485[1]; // @[OneHot.scala 66:30:@41008.4]
  assign _T_96488 = _T_96485[2]; // @[OneHot.scala 66:30:@41009.4]
  assign _T_96489 = _T_96485[3]; // @[OneHot.scala 66:30:@41010.4]
  assign _T_96490 = _T_96485[4]; // @[OneHot.scala 66:30:@41011.4]
  assign _T_96491 = _T_96485[5]; // @[OneHot.scala 66:30:@41012.4]
  assign _T_96492 = _T_96485[6]; // @[OneHot.scala 66:30:@41013.4]
  assign _T_96493 = _T_96485[7]; // @[OneHot.scala 66:30:@41014.4]
  assign _T_96494 = _T_96485[8]; // @[OneHot.scala 66:30:@41015.4]
  assign _T_96495 = _T_96485[9]; // @[OneHot.scala 66:30:@41016.4]
  assign _T_96496 = _T_96485[10]; // @[OneHot.scala 66:30:@41017.4]
  assign _T_96497 = _T_96485[11]; // @[OneHot.scala 66:30:@41018.4]
  assign _T_96498 = _T_96485[12]; // @[OneHot.scala 66:30:@41019.4]
  assign _T_96499 = _T_96485[13]; // @[OneHot.scala 66:30:@41020.4]
  assign _T_96500 = _T_96485[14]; // @[OneHot.scala 66:30:@41021.4]
  assign _T_96501 = _T_96485[15]; // @[OneHot.scala 66:30:@41022.4]
  assign _T_96542 = entriesPorts_0_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41040.4]
  assign _T_96543 = entriesPorts_0_6 ? 16'h4000 : _T_96542; // @[Mux.scala 31:69:@41041.4]
  assign _T_96544 = entriesPorts_0_5 ? 16'h2000 : _T_96543; // @[Mux.scala 31:69:@41042.4]
  assign _T_96545 = entriesPorts_0_4 ? 16'h1000 : _T_96544; // @[Mux.scala 31:69:@41043.4]
  assign _T_96546 = entriesPorts_0_3 ? 16'h800 : _T_96545; // @[Mux.scala 31:69:@41044.4]
  assign _T_96547 = entriesPorts_0_2 ? 16'h400 : _T_96546; // @[Mux.scala 31:69:@41045.4]
  assign _T_96548 = entriesPorts_0_1 ? 16'h200 : _T_96547; // @[Mux.scala 31:69:@41046.4]
  assign _T_96549 = entriesPorts_0_0 ? 16'h100 : _T_96548; // @[Mux.scala 31:69:@41047.4]
  assign _T_96550 = entriesPorts_0_15 ? 16'h80 : _T_96549; // @[Mux.scala 31:69:@41048.4]
  assign _T_96551 = entriesPorts_0_14 ? 16'h40 : _T_96550; // @[Mux.scala 31:69:@41049.4]
  assign _T_96552 = entriesPorts_0_13 ? 16'h20 : _T_96551; // @[Mux.scala 31:69:@41050.4]
  assign _T_96553 = entriesPorts_0_12 ? 16'h10 : _T_96552; // @[Mux.scala 31:69:@41051.4]
  assign _T_96554 = entriesPorts_0_11 ? 16'h8 : _T_96553; // @[Mux.scala 31:69:@41052.4]
  assign _T_96555 = entriesPorts_0_10 ? 16'h4 : _T_96554; // @[Mux.scala 31:69:@41053.4]
  assign _T_96556 = entriesPorts_0_9 ? 16'h2 : _T_96555; // @[Mux.scala 31:69:@41054.4]
  assign _T_96557 = entriesPorts_0_8 ? 16'h1 : _T_96556; // @[Mux.scala 31:69:@41055.4]
  assign _T_96558 = _T_96557[0]; // @[OneHot.scala 66:30:@41056.4]
  assign _T_96559 = _T_96557[1]; // @[OneHot.scala 66:30:@41057.4]
  assign _T_96560 = _T_96557[2]; // @[OneHot.scala 66:30:@41058.4]
  assign _T_96561 = _T_96557[3]; // @[OneHot.scala 66:30:@41059.4]
  assign _T_96562 = _T_96557[4]; // @[OneHot.scala 66:30:@41060.4]
  assign _T_96563 = _T_96557[5]; // @[OneHot.scala 66:30:@41061.4]
  assign _T_96564 = _T_96557[6]; // @[OneHot.scala 66:30:@41062.4]
  assign _T_96565 = _T_96557[7]; // @[OneHot.scala 66:30:@41063.4]
  assign _T_96566 = _T_96557[8]; // @[OneHot.scala 66:30:@41064.4]
  assign _T_96567 = _T_96557[9]; // @[OneHot.scala 66:30:@41065.4]
  assign _T_96568 = _T_96557[10]; // @[OneHot.scala 66:30:@41066.4]
  assign _T_96569 = _T_96557[11]; // @[OneHot.scala 66:30:@41067.4]
  assign _T_96570 = _T_96557[12]; // @[OneHot.scala 66:30:@41068.4]
  assign _T_96571 = _T_96557[13]; // @[OneHot.scala 66:30:@41069.4]
  assign _T_96572 = _T_96557[14]; // @[OneHot.scala 66:30:@41070.4]
  assign _T_96573 = _T_96557[15]; // @[OneHot.scala 66:30:@41071.4]
  assign _T_96614 = entriesPorts_0_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41089.4]
  assign _T_96615 = entriesPorts_0_7 ? 16'h4000 : _T_96614; // @[Mux.scala 31:69:@41090.4]
  assign _T_96616 = entriesPorts_0_6 ? 16'h2000 : _T_96615; // @[Mux.scala 31:69:@41091.4]
  assign _T_96617 = entriesPorts_0_5 ? 16'h1000 : _T_96616; // @[Mux.scala 31:69:@41092.4]
  assign _T_96618 = entriesPorts_0_4 ? 16'h800 : _T_96617; // @[Mux.scala 31:69:@41093.4]
  assign _T_96619 = entriesPorts_0_3 ? 16'h400 : _T_96618; // @[Mux.scala 31:69:@41094.4]
  assign _T_96620 = entriesPorts_0_2 ? 16'h200 : _T_96619; // @[Mux.scala 31:69:@41095.4]
  assign _T_96621 = entriesPorts_0_1 ? 16'h100 : _T_96620; // @[Mux.scala 31:69:@41096.4]
  assign _T_96622 = entriesPorts_0_0 ? 16'h80 : _T_96621; // @[Mux.scala 31:69:@41097.4]
  assign _T_96623 = entriesPorts_0_15 ? 16'h40 : _T_96622; // @[Mux.scala 31:69:@41098.4]
  assign _T_96624 = entriesPorts_0_14 ? 16'h20 : _T_96623; // @[Mux.scala 31:69:@41099.4]
  assign _T_96625 = entriesPorts_0_13 ? 16'h10 : _T_96624; // @[Mux.scala 31:69:@41100.4]
  assign _T_96626 = entriesPorts_0_12 ? 16'h8 : _T_96625; // @[Mux.scala 31:69:@41101.4]
  assign _T_96627 = entriesPorts_0_11 ? 16'h4 : _T_96626; // @[Mux.scala 31:69:@41102.4]
  assign _T_96628 = entriesPorts_0_10 ? 16'h2 : _T_96627; // @[Mux.scala 31:69:@41103.4]
  assign _T_96629 = entriesPorts_0_9 ? 16'h1 : _T_96628; // @[Mux.scala 31:69:@41104.4]
  assign _T_96630 = _T_96629[0]; // @[OneHot.scala 66:30:@41105.4]
  assign _T_96631 = _T_96629[1]; // @[OneHot.scala 66:30:@41106.4]
  assign _T_96632 = _T_96629[2]; // @[OneHot.scala 66:30:@41107.4]
  assign _T_96633 = _T_96629[3]; // @[OneHot.scala 66:30:@41108.4]
  assign _T_96634 = _T_96629[4]; // @[OneHot.scala 66:30:@41109.4]
  assign _T_96635 = _T_96629[5]; // @[OneHot.scala 66:30:@41110.4]
  assign _T_96636 = _T_96629[6]; // @[OneHot.scala 66:30:@41111.4]
  assign _T_96637 = _T_96629[7]; // @[OneHot.scala 66:30:@41112.4]
  assign _T_96638 = _T_96629[8]; // @[OneHot.scala 66:30:@41113.4]
  assign _T_96639 = _T_96629[9]; // @[OneHot.scala 66:30:@41114.4]
  assign _T_96640 = _T_96629[10]; // @[OneHot.scala 66:30:@41115.4]
  assign _T_96641 = _T_96629[11]; // @[OneHot.scala 66:30:@41116.4]
  assign _T_96642 = _T_96629[12]; // @[OneHot.scala 66:30:@41117.4]
  assign _T_96643 = _T_96629[13]; // @[OneHot.scala 66:30:@41118.4]
  assign _T_96644 = _T_96629[14]; // @[OneHot.scala 66:30:@41119.4]
  assign _T_96645 = _T_96629[15]; // @[OneHot.scala 66:30:@41120.4]
  assign _T_96686 = entriesPorts_0_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41138.4]
  assign _T_96687 = entriesPorts_0_8 ? 16'h4000 : _T_96686; // @[Mux.scala 31:69:@41139.4]
  assign _T_96688 = entriesPorts_0_7 ? 16'h2000 : _T_96687; // @[Mux.scala 31:69:@41140.4]
  assign _T_96689 = entriesPorts_0_6 ? 16'h1000 : _T_96688; // @[Mux.scala 31:69:@41141.4]
  assign _T_96690 = entriesPorts_0_5 ? 16'h800 : _T_96689; // @[Mux.scala 31:69:@41142.4]
  assign _T_96691 = entriesPorts_0_4 ? 16'h400 : _T_96690; // @[Mux.scala 31:69:@41143.4]
  assign _T_96692 = entriesPorts_0_3 ? 16'h200 : _T_96691; // @[Mux.scala 31:69:@41144.4]
  assign _T_96693 = entriesPorts_0_2 ? 16'h100 : _T_96692; // @[Mux.scala 31:69:@41145.4]
  assign _T_96694 = entriesPorts_0_1 ? 16'h80 : _T_96693; // @[Mux.scala 31:69:@41146.4]
  assign _T_96695 = entriesPorts_0_0 ? 16'h40 : _T_96694; // @[Mux.scala 31:69:@41147.4]
  assign _T_96696 = entriesPorts_0_15 ? 16'h20 : _T_96695; // @[Mux.scala 31:69:@41148.4]
  assign _T_96697 = entriesPorts_0_14 ? 16'h10 : _T_96696; // @[Mux.scala 31:69:@41149.4]
  assign _T_96698 = entriesPorts_0_13 ? 16'h8 : _T_96697; // @[Mux.scala 31:69:@41150.4]
  assign _T_96699 = entriesPorts_0_12 ? 16'h4 : _T_96698; // @[Mux.scala 31:69:@41151.4]
  assign _T_96700 = entriesPorts_0_11 ? 16'h2 : _T_96699; // @[Mux.scala 31:69:@41152.4]
  assign _T_96701 = entriesPorts_0_10 ? 16'h1 : _T_96700; // @[Mux.scala 31:69:@41153.4]
  assign _T_96702 = _T_96701[0]; // @[OneHot.scala 66:30:@41154.4]
  assign _T_96703 = _T_96701[1]; // @[OneHot.scala 66:30:@41155.4]
  assign _T_96704 = _T_96701[2]; // @[OneHot.scala 66:30:@41156.4]
  assign _T_96705 = _T_96701[3]; // @[OneHot.scala 66:30:@41157.4]
  assign _T_96706 = _T_96701[4]; // @[OneHot.scala 66:30:@41158.4]
  assign _T_96707 = _T_96701[5]; // @[OneHot.scala 66:30:@41159.4]
  assign _T_96708 = _T_96701[6]; // @[OneHot.scala 66:30:@41160.4]
  assign _T_96709 = _T_96701[7]; // @[OneHot.scala 66:30:@41161.4]
  assign _T_96710 = _T_96701[8]; // @[OneHot.scala 66:30:@41162.4]
  assign _T_96711 = _T_96701[9]; // @[OneHot.scala 66:30:@41163.4]
  assign _T_96712 = _T_96701[10]; // @[OneHot.scala 66:30:@41164.4]
  assign _T_96713 = _T_96701[11]; // @[OneHot.scala 66:30:@41165.4]
  assign _T_96714 = _T_96701[12]; // @[OneHot.scala 66:30:@41166.4]
  assign _T_96715 = _T_96701[13]; // @[OneHot.scala 66:30:@41167.4]
  assign _T_96716 = _T_96701[14]; // @[OneHot.scala 66:30:@41168.4]
  assign _T_96717 = _T_96701[15]; // @[OneHot.scala 66:30:@41169.4]
  assign _T_96758 = entriesPorts_0_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41187.4]
  assign _T_96759 = entriesPorts_0_9 ? 16'h4000 : _T_96758; // @[Mux.scala 31:69:@41188.4]
  assign _T_96760 = entriesPorts_0_8 ? 16'h2000 : _T_96759; // @[Mux.scala 31:69:@41189.4]
  assign _T_96761 = entriesPorts_0_7 ? 16'h1000 : _T_96760; // @[Mux.scala 31:69:@41190.4]
  assign _T_96762 = entriesPorts_0_6 ? 16'h800 : _T_96761; // @[Mux.scala 31:69:@41191.4]
  assign _T_96763 = entriesPorts_0_5 ? 16'h400 : _T_96762; // @[Mux.scala 31:69:@41192.4]
  assign _T_96764 = entriesPorts_0_4 ? 16'h200 : _T_96763; // @[Mux.scala 31:69:@41193.4]
  assign _T_96765 = entriesPorts_0_3 ? 16'h100 : _T_96764; // @[Mux.scala 31:69:@41194.4]
  assign _T_96766 = entriesPorts_0_2 ? 16'h80 : _T_96765; // @[Mux.scala 31:69:@41195.4]
  assign _T_96767 = entriesPorts_0_1 ? 16'h40 : _T_96766; // @[Mux.scala 31:69:@41196.4]
  assign _T_96768 = entriesPorts_0_0 ? 16'h20 : _T_96767; // @[Mux.scala 31:69:@41197.4]
  assign _T_96769 = entriesPorts_0_15 ? 16'h10 : _T_96768; // @[Mux.scala 31:69:@41198.4]
  assign _T_96770 = entriesPorts_0_14 ? 16'h8 : _T_96769; // @[Mux.scala 31:69:@41199.4]
  assign _T_96771 = entriesPorts_0_13 ? 16'h4 : _T_96770; // @[Mux.scala 31:69:@41200.4]
  assign _T_96772 = entriesPorts_0_12 ? 16'h2 : _T_96771; // @[Mux.scala 31:69:@41201.4]
  assign _T_96773 = entriesPorts_0_11 ? 16'h1 : _T_96772; // @[Mux.scala 31:69:@41202.4]
  assign _T_96774 = _T_96773[0]; // @[OneHot.scala 66:30:@41203.4]
  assign _T_96775 = _T_96773[1]; // @[OneHot.scala 66:30:@41204.4]
  assign _T_96776 = _T_96773[2]; // @[OneHot.scala 66:30:@41205.4]
  assign _T_96777 = _T_96773[3]; // @[OneHot.scala 66:30:@41206.4]
  assign _T_96778 = _T_96773[4]; // @[OneHot.scala 66:30:@41207.4]
  assign _T_96779 = _T_96773[5]; // @[OneHot.scala 66:30:@41208.4]
  assign _T_96780 = _T_96773[6]; // @[OneHot.scala 66:30:@41209.4]
  assign _T_96781 = _T_96773[7]; // @[OneHot.scala 66:30:@41210.4]
  assign _T_96782 = _T_96773[8]; // @[OneHot.scala 66:30:@41211.4]
  assign _T_96783 = _T_96773[9]; // @[OneHot.scala 66:30:@41212.4]
  assign _T_96784 = _T_96773[10]; // @[OneHot.scala 66:30:@41213.4]
  assign _T_96785 = _T_96773[11]; // @[OneHot.scala 66:30:@41214.4]
  assign _T_96786 = _T_96773[12]; // @[OneHot.scala 66:30:@41215.4]
  assign _T_96787 = _T_96773[13]; // @[OneHot.scala 66:30:@41216.4]
  assign _T_96788 = _T_96773[14]; // @[OneHot.scala 66:30:@41217.4]
  assign _T_96789 = _T_96773[15]; // @[OneHot.scala 66:30:@41218.4]
  assign _T_96830 = entriesPorts_0_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41236.4]
  assign _T_96831 = entriesPorts_0_10 ? 16'h4000 : _T_96830; // @[Mux.scala 31:69:@41237.4]
  assign _T_96832 = entriesPorts_0_9 ? 16'h2000 : _T_96831; // @[Mux.scala 31:69:@41238.4]
  assign _T_96833 = entriesPorts_0_8 ? 16'h1000 : _T_96832; // @[Mux.scala 31:69:@41239.4]
  assign _T_96834 = entriesPorts_0_7 ? 16'h800 : _T_96833; // @[Mux.scala 31:69:@41240.4]
  assign _T_96835 = entriesPorts_0_6 ? 16'h400 : _T_96834; // @[Mux.scala 31:69:@41241.4]
  assign _T_96836 = entriesPorts_0_5 ? 16'h200 : _T_96835; // @[Mux.scala 31:69:@41242.4]
  assign _T_96837 = entriesPorts_0_4 ? 16'h100 : _T_96836; // @[Mux.scala 31:69:@41243.4]
  assign _T_96838 = entriesPorts_0_3 ? 16'h80 : _T_96837; // @[Mux.scala 31:69:@41244.4]
  assign _T_96839 = entriesPorts_0_2 ? 16'h40 : _T_96838; // @[Mux.scala 31:69:@41245.4]
  assign _T_96840 = entriesPorts_0_1 ? 16'h20 : _T_96839; // @[Mux.scala 31:69:@41246.4]
  assign _T_96841 = entriesPorts_0_0 ? 16'h10 : _T_96840; // @[Mux.scala 31:69:@41247.4]
  assign _T_96842 = entriesPorts_0_15 ? 16'h8 : _T_96841; // @[Mux.scala 31:69:@41248.4]
  assign _T_96843 = entriesPorts_0_14 ? 16'h4 : _T_96842; // @[Mux.scala 31:69:@41249.4]
  assign _T_96844 = entriesPorts_0_13 ? 16'h2 : _T_96843; // @[Mux.scala 31:69:@41250.4]
  assign _T_96845 = entriesPorts_0_12 ? 16'h1 : _T_96844; // @[Mux.scala 31:69:@41251.4]
  assign _T_96846 = _T_96845[0]; // @[OneHot.scala 66:30:@41252.4]
  assign _T_96847 = _T_96845[1]; // @[OneHot.scala 66:30:@41253.4]
  assign _T_96848 = _T_96845[2]; // @[OneHot.scala 66:30:@41254.4]
  assign _T_96849 = _T_96845[3]; // @[OneHot.scala 66:30:@41255.4]
  assign _T_96850 = _T_96845[4]; // @[OneHot.scala 66:30:@41256.4]
  assign _T_96851 = _T_96845[5]; // @[OneHot.scala 66:30:@41257.4]
  assign _T_96852 = _T_96845[6]; // @[OneHot.scala 66:30:@41258.4]
  assign _T_96853 = _T_96845[7]; // @[OneHot.scala 66:30:@41259.4]
  assign _T_96854 = _T_96845[8]; // @[OneHot.scala 66:30:@41260.4]
  assign _T_96855 = _T_96845[9]; // @[OneHot.scala 66:30:@41261.4]
  assign _T_96856 = _T_96845[10]; // @[OneHot.scala 66:30:@41262.4]
  assign _T_96857 = _T_96845[11]; // @[OneHot.scala 66:30:@41263.4]
  assign _T_96858 = _T_96845[12]; // @[OneHot.scala 66:30:@41264.4]
  assign _T_96859 = _T_96845[13]; // @[OneHot.scala 66:30:@41265.4]
  assign _T_96860 = _T_96845[14]; // @[OneHot.scala 66:30:@41266.4]
  assign _T_96861 = _T_96845[15]; // @[OneHot.scala 66:30:@41267.4]
  assign _T_96902 = entriesPorts_0_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41285.4]
  assign _T_96903 = entriesPorts_0_11 ? 16'h4000 : _T_96902; // @[Mux.scala 31:69:@41286.4]
  assign _T_96904 = entriesPorts_0_10 ? 16'h2000 : _T_96903; // @[Mux.scala 31:69:@41287.4]
  assign _T_96905 = entriesPorts_0_9 ? 16'h1000 : _T_96904; // @[Mux.scala 31:69:@41288.4]
  assign _T_96906 = entriesPorts_0_8 ? 16'h800 : _T_96905; // @[Mux.scala 31:69:@41289.4]
  assign _T_96907 = entriesPorts_0_7 ? 16'h400 : _T_96906; // @[Mux.scala 31:69:@41290.4]
  assign _T_96908 = entriesPorts_0_6 ? 16'h200 : _T_96907; // @[Mux.scala 31:69:@41291.4]
  assign _T_96909 = entriesPorts_0_5 ? 16'h100 : _T_96908; // @[Mux.scala 31:69:@41292.4]
  assign _T_96910 = entriesPorts_0_4 ? 16'h80 : _T_96909; // @[Mux.scala 31:69:@41293.4]
  assign _T_96911 = entriesPorts_0_3 ? 16'h40 : _T_96910; // @[Mux.scala 31:69:@41294.4]
  assign _T_96912 = entriesPorts_0_2 ? 16'h20 : _T_96911; // @[Mux.scala 31:69:@41295.4]
  assign _T_96913 = entriesPorts_0_1 ? 16'h10 : _T_96912; // @[Mux.scala 31:69:@41296.4]
  assign _T_96914 = entriesPorts_0_0 ? 16'h8 : _T_96913; // @[Mux.scala 31:69:@41297.4]
  assign _T_96915 = entriesPorts_0_15 ? 16'h4 : _T_96914; // @[Mux.scala 31:69:@41298.4]
  assign _T_96916 = entriesPorts_0_14 ? 16'h2 : _T_96915; // @[Mux.scala 31:69:@41299.4]
  assign _T_96917 = entriesPorts_0_13 ? 16'h1 : _T_96916; // @[Mux.scala 31:69:@41300.4]
  assign _T_96918 = _T_96917[0]; // @[OneHot.scala 66:30:@41301.4]
  assign _T_96919 = _T_96917[1]; // @[OneHot.scala 66:30:@41302.4]
  assign _T_96920 = _T_96917[2]; // @[OneHot.scala 66:30:@41303.4]
  assign _T_96921 = _T_96917[3]; // @[OneHot.scala 66:30:@41304.4]
  assign _T_96922 = _T_96917[4]; // @[OneHot.scala 66:30:@41305.4]
  assign _T_96923 = _T_96917[5]; // @[OneHot.scala 66:30:@41306.4]
  assign _T_96924 = _T_96917[6]; // @[OneHot.scala 66:30:@41307.4]
  assign _T_96925 = _T_96917[7]; // @[OneHot.scala 66:30:@41308.4]
  assign _T_96926 = _T_96917[8]; // @[OneHot.scala 66:30:@41309.4]
  assign _T_96927 = _T_96917[9]; // @[OneHot.scala 66:30:@41310.4]
  assign _T_96928 = _T_96917[10]; // @[OneHot.scala 66:30:@41311.4]
  assign _T_96929 = _T_96917[11]; // @[OneHot.scala 66:30:@41312.4]
  assign _T_96930 = _T_96917[12]; // @[OneHot.scala 66:30:@41313.4]
  assign _T_96931 = _T_96917[13]; // @[OneHot.scala 66:30:@41314.4]
  assign _T_96932 = _T_96917[14]; // @[OneHot.scala 66:30:@41315.4]
  assign _T_96933 = _T_96917[15]; // @[OneHot.scala 66:30:@41316.4]
  assign _T_96974 = entriesPorts_0_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41334.4]
  assign _T_96975 = entriesPorts_0_12 ? 16'h4000 : _T_96974; // @[Mux.scala 31:69:@41335.4]
  assign _T_96976 = entriesPorts_0_11 ? 16'h2000 : _T_96975; // @[Mux.scala 31:69:@41336.4]
  assign _T_96977 = entriesPorts_0_10 ? 16'h1000 : _T_96976; // @[Mux.scala 31:69:@41337.4]
  assign _T_96978 = entriesPorts_0_9 ? 16'h800 : _T_96977; // @[Mux.scala 31:69:@41338.4]
  assign _T_96979 = entriesPorts_0_8 ? 16'h400 : _T_96978; // @[Mux.scala 31:69:@41339.4]
  assign _T_96980 = entriesPorts_0_7 ? 16'h200 : _T_96979; // @[Mux.scala 31:69:@41340.4]
  assign _T_96981 = entriesPorts_0_6 ? 16'h100 : _T_96980; // @[Mux.scala 31:69:@41341.4]
  assign _T_96982 = entriesPorts_0_5 ? 16'h80 : _T_96981; // @[Mux.scala 31:69:@41342.4]
  assign _T_96983 = entriesPorts_0_4 ? 16'h40 : _T_96982; // @[Mux.scala 31:69:@41343.4]
  assign _T_96984 = entriesPorts_0_3 ? 16'h20 : _T_96983; // @[Mux.scala 31:69:@41344.4]
  assign _T_96985 = entriesPorts_0_2 ? 16'h10 : _T_96984; // @[Mux.scala 31:69:@41345.4]
  assign _T_96986 = entriesPorts_0_1 ? 16'h8 : _T_96985; // @[Mux.scala 31:69:@41346.4]
  assign _T_96987 = entriesPorts_0_0 ? 16'h4 : _T_96986; // @[Mux.scala 31:69:@41347.4]
  assign _T_96988 = entriesPorts_0_15 ? 16'h2 : _T_96987; // @[Mux.scala 31:69:@41348.4]
  assign _T_96989 = entriesPorts_0_14 ? 16'h1 : _T_96988; // @[Mux.scala 31:69:@41349.4]
  assign _T_96990 = _T_96989[0]; // @[OneHot.scala 66:30:@41350.4]
  assign _T_96991 = _T_96989[1]; // @[OneHot.scala 66:30:@41351.4]
  assign _T_96992 = _T_96989[2]; // @[OneHot.scala 66:30:@41352.4]
  assign _T_96993 = _T_96989[3]; // @[OneHot.scala 66:30:@41353.4]
  assign _T_96994 = _T_96989[4]; // @[OneHot.scala 66:30:@41354.4]
  assign _T_96995 = _T_96989[5]; // @[OneHot.scala 66:30:@41355.4]
  assign _T_96996 = _T_96989[6]; // @[OneHot.scala 66:30:@41356.4]
  assign _T_96997 = _T_96989[7]; // @[OneHot.scala 66:30:@41357.4]
  assign _T_96998 = _T_96989[8]; // @[OneHot.scala 66:30:@41358.4]
  assign _T_96999 = _T_96989[9]; // @[OneHot.scala 66:30:@41359.4]
  assign _T_97000 = _T_96989[10]; // @[OneHot.scala 66:30:@41360.4]
  assign _T_97001 = _T_96989[11]; // @[OneHot.scala 66:30:@41361.4]
  assign _T_97002 = _T_96989[12]; // @[OneHot.scala 66:30:@41362.4]
  assign _T_97003 = _T_96989[13]; // @[OneHot.scala 66:30:@41363.4]
  assign _T_97004 = _T_96989[14]; // @[OneHot.scala 66:30:@41364.4]
  assign _T_97005 = _T_96989[15]; // @[OneHot.scala 66:30:@41365.4]
  assign _T_97046 = entriesPorts_0_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41383.4]
  assign _T_97047 = entriesPorts_0_13 ? 16'h4000 : _T_97046; // @[Mux.scala 31:69:@41384.4]
  assign _T_97048 = entriesPorts_0_12 ? 16'h2000 : _T_97047; // @[Mux.scala 31:69:@41385.4]
  assign _T_97049 = entriesPorts_0_11 ? 16'h1000 : _T_97048; // @[Mux.scala 31:69:@41386.4]
  assign _T_97050 = entriesPorts_0_10 ? 16'h800 : _T_97049; // @[Mux.scala 31:69:@41387.4]
  assign _T_97051 = entriesPorts_0_9 ? 16'h400 : _T_97050; // @[Mux.scala 31:69:@41388.4]
  assign _T_97052 = entriesPorts_0_8 ? 16'h200 : _T_97051; // @[Mux.scala 31:69:@41389.4]
  assign _T_97053 = entriesPorts_0_7 ? 16'h100 : _T_97052; // @[Mux.scala 31:69:@41390.4]
  assign _T_97054 = entriesPorts_0_6 ? 16'h80 : _T_97053; // @[Mux.scala 31:69:@41391.4]
  assign _T_97055 = entriesPorts_0_5 ? 16'h40 : _T_97054; // @[Mux.scala 31:69:@41392.4]
  assign _T_97056 = entriesPorts_0_4 ? 16'h20 : _T_97055; // @[Mux.scala 31:69:@41393.4]
  assign _T_97057 = entriesPorts_0_3 ? 16'h10 : _T_97056; // @[Mux.scala 31:69:@41394.4]
  assign _T_97058 = entriesPorts_0_2 ? 16'h8 : _T_97057; // @[Mux.scala 31:69:@41395.4]
  assign _T_97059 = entriesPorts_0_1 ? 16'h4 : _T_97058; // @[Mux.scala 31:69:@41396.4]
  assign _T_97060 = entriesPorts_0_0 ? 16'h2 : _T_97059; // @[Mux.scala 31:69:@41397.4]
  assign _T_97061 = entriesPorts_0_15 ? 16'h1 : _T_97060; // @[Mux.scala 31:69:@41398.4]
  assign _T_97062 = _T_97061[0]; // @[OneHot.scala 66:30:@41399.4]
  assign _T_97063 = _T_97061[1]; // @[OneHot.scala 66:30:@41400.4]
  assign _T_97064 = _T_97061[2]; // @[OneHot.scala 66:30:@41401.4]
  assign _T_97065 = _T_97061[3]; // @[OneHot.scala 66:30:@41402.4]
  assign _T_97066 = _T_97061[4]; // @[OneHot.scala 66:30:@41403.4]
  assign _T_97067 = _T_97061[5]; // @[OneHot.scala 66:30:@41404.4]
  assign _T_97068 = _T_97061[6]; // @[OneHot.scala 66:30:@41405.4]
  assign _T_97069 = _T_97061[7]; // @[OneHot.scala 66:30:@41406.4]
  assign _T_97070 = _T_97061[8]; // @[OneHot.scala 66:30:@41407.4]
  assign _T_97071 = _T_97061[9]; // @[OneHot.scala 66:30:@41408.4]
  assign _T_97072 = _T_97061[10]; // @[OneHot.scala 66:30:@41409.4]
  assign _T_97073 = _T_97061[11]; // @[OneHot.scala 66:30:@41410.4]
  assign _T_97074 = _T_97061[12]; // @[OneHot.scala 66:30:@41411.4]
  assign _T_97075 = _T_97061[13]; // @[OneHot.scala 66:30:@41412.4]
  assign _T_97076 = _T_97061[14]; // @[OneHot.scala 66:30:@41413.4]
  assign _T_97077 = _T_97061[15]; // @[OneHot.scala 66:30:@41414.4]
  assign _T_97142 = {_T_95989,_T_95988,_T_95987,_T_95986,_T_95985,_T_95984,_T_95983,_T_95982}; // @[Mux.scala 19:72:@41438.4]
  assign _T_97150 = {_T_95997,_T_95996,_T_95995,_T_95994,_T_95993,_T_95992,_T_95991,_T_95990,_T_97142}; // @[Mux.scala 19:72:@41446.4]
  assign _T_97152 = _T_90400 ? _T_97150 : 16'h0; // @[Mux.scala 19:72:@41447.4]
  assign _T_97159 = {_T_96060,_T_96059,_T_96058,_T_96057,_T_96056,_T_96055,_T_96054,_T_96069}; // @[Mux.scala 19:72:@41454.4]
  assign _T_97167 = {_T_96068,_T_96067,_T_96066,_T_96065,_T_96064,_T_96063,_T_96062,_T_96061,_T_97159}; // @[Mux.scala 19:72:@41462.4]
  assign _T_97169 = _T_90401 ? _T_97167 : 16'h0; // @[Mux.scala 19:72:@41463.4]
  assign _T_97176 = {_T_96131,_T_96130,_T_96129,_T_96128,_T_96127,_T_96126,_T_96141,_T_96140}; // @[Mux.scala 19:72:@41470.4]
  assign _T_97184 = {_T_96139,_T_96138,_T_96137,_T_96136,_T_96135,_T_96134,_T_96133,_T_96132,_T_97176}; // @[Mux.scala 19:72:@41478.4]
  assign _T_97186 = _T_90402 ? _T_97184 : 16'h0; // @[Mux.scala 19:72:@41479.4]
  assign _T_97193 = {_T_96202,_T_96201,_T_96200,_T_96199,_T_96198,_T_96213,_T_96212,_T_96211}; // @[Mux.scala 19:72:@41486.4]
  assign _T_97201 = {_T_96210,_T_96209,_T_96208,_T_96207,_T_96206,_T_96205,_T_96204,_T_96203,_T_97193}; // @[Mux.scala 19:72:@41494.4]
  assign _T_97203 = _T_90403 ? _T_97201 : 16'h0; // @[Mux.scala 19:72:@41495.4]
  assign _T_97210 = {_T_96273,_T_96272,_T_96271,_T_96270,_T_96285,_T_96284,_T_96283,_T_96282}; // @[Mux.scala 19:72:@41502.4]
  assign _T_97218 = {_T_96281,_T_96280,_T_96279,_T_96278,_T_96277,_T_96276,_T_96275,_T_96274,_T_97210}; // @[Mux.scala 19:72:@41510.4]
  assign _T_97220 = _T_90404 ? _T_97218 : 16'h0; // @[Mux.scala 19:72:@41511.4]
  assign _T_97227 = {_T_96344,_T_96343,_T_96342,_T_96357,_T_96356,_T_96355,_T_96354,_T_96353}; // @[Mux.scala 19:72:@41518.4]
  assign _T_97235 = {_T_96352,_T_96351,_T_96350,_T_96349,_T_96348,_T_96347,_T_96346,_T_96345,_T_97227}; // @[Mux.scala 19:72:@41526.4]
  assign _T_97237 = _T_90405 ? _T_97235 : 16'h0; // @[Mux.scala 19:72:@41527.4]
  assign _T_97244 = {_T_96415,_T_96414,_T_96429,_T_96428,_T_96427,_T_96426,_T_96425,_T_96424}; // @[Mux.scala 19:72:@41534.4]
  assign _T_97252 = {_T_96423,_T_96422,_T_96421,_T_96420,_T_96419,_T_96418,_T_96417,_T_96416,_T_97244}; // @[Mux.scala 19:72:@41542.4]
  assign _T_97254 = _T_90406 ? _T_97252 : 16'h0; // @[Mux.scala 19:72:@41543.4]
  assign _T_97261 = {_T_96486,_T_96501,_T_96500,_T_96499,_T_96498,_T_96497,_T_96496,_T_96495}; // @[Mux.scala 19:72:@41550.4]
  assign _T_97269 = {_T_96494,_T_96493,_T_96492,_T_96491,_T_96490,_T_96489,_T_96488,_T_96487,_T_97261}; // @[Mux.scala 19:72:@41558.4]
  assign _T_97271 = _T_90407 ? _T_97269 : 16'h0; // @[Mux.scala 19:72:@41559.4]
  assign _T_97278 = {_T_96573,_T_96572,_T_96571,_T_96570,_T_96569,_T_96568,_T_96567,_T_96566}; // @[Mux.scala 19:72:@41566.4]
  assign _T_97286 = {_T_96565,_T_96564,_T_96563,_T_96562,_T_96561,_T_96560,_T_96559,_T_96558,_T_97278}; // @[Mux.scala 19:72:@41574.4]
  assign _T_97288 = _T_90408 ? _T_97286 : 16'h0; // @[Mux.scala 19:72:@41575.4]
  assign _T_97295 = {_T_96644,_T_96643,_T_96642,_T_96641,_T_96640,_T_96639,_T_96638,_T_96637}; // @[Mux.scala 19:72:@41582.4]
  assign _T_97303 = {_T_96636,_T_96635,_T_96634,_T_96633,_T_96632,_T_96631,_T_96630,_T_96645,_T_97295}; // @[Mux.scala 19:72:@41590.4]
  assign _T_97305 = _T_90409 ? _T_97303 : 16'h0; // @[Mux.scala 19:72:@41591.4]
  assign _T_97312 = {_T_96715,_T_96714,_T_96713,_T_96712,_T_96711,_T_96710,_T_96709,_T_96708}; // @[Mux.scala 19:72:@41598.4]
  assign _T_97320 = {_T_96707,_T_96706,_T_96705,_T_96704,_T_96703,_T_96702,_T_96717,_T_96716,_T_97312}; // @[Mux.scala 19:72:@41606.4]
  assign _T_97322 = _T_90410 ? _T_97320 : 16'h0; // @[Mux.scala 19:72:@41607.4]
  assign _T_97329 = {_T_96786,_T_96785,_T_96784,_T_96783,_T_96782,_T_96781,_T_96780,_T_96779}; // @[Mux.scala 19:72:@41614.4]
  assign _T_97337 = {_T_96778,_T_96777,_T_96776,_T_96775,_T_96774,_T_96789,_T_96788,_T_96787,_T_97329}; // @[Mux.scala 19:72:@41622.4]
  assign _T_97339 = _T_90411 ? _T_97337 : 16'h0; // @[Mux.scala 19:72:@41623.4]
  assign _T_97346 = {_T_96857,_T_96856,_T_96855,_T_96854,_T_96853,_T_96852,_T_96851,_T_96850}; // @[Mux.scala 19:72:@41630.4]
  assign _T_97354 = {_T_96849,_T_96848,_T_96847,_T_96846,_T_96861,_T_96860,_T_96859,_T_96858,_T_97346}; // @[Mux.scala 19:72:@41638.4]
  assign _T_97356 = _T_90412 ? _T_97354 : 16'h0; // @[Mux.scala 19:72:@41639.4]
  assign _T_97363 = {_T_96928,_T_96927,_T_96926,_T_96925,_T_96924,_T_96923,_T_96922,_T_96921}; // @[Mux.scala 19:72:@41646.4]
  assign _T_97371 = {_T_96920,_T_96919,_T_96918,_T_96933,_T_96932,_T_96931,_T_96930,_T_96929,_T_97363}; // @[Mux.scala 19:72:@41654.4]
  assign _T_97373 = _T_90413 ? _T_97371 : 16'h0; // @[Mux.scala 19:72:@41655.4]
  assign _T_97380 = {_T_96999,_T_96998,_T_96997,_T_96996,_T_96995,_T_96994,_T_96993,_T_96992}; // @[Mux.scala 19:72:@41662.4]
  assign _T_97388 = {_T_96991,_T_96990,_T_97005,_T_97004,_T_97003,_T_97002,_T_97001,_T_97000,_T_97380}; // @[Mux.scala 19:72:@41670.4]
  assign _T_97390 = _T_90414 ? _T_97388 : 16'h0; // @[Mux.scala 19:72:@41671.4]
  assign _T_97397 = {_T_97070,_T_97069,_T_97068,_T_97067,_T_97066,_T_97065,_T_97064,_T_97063}; // @[Mux.scala 19:72:@41678.4]
  assign _T_97405 = {_T_97062,_T_97077,_T_97076,_T_97075,_T_97074,_T_97073,_T_97072,_T_97071,_T_97397}; // @[Mux.scala 19:72:@41686.4]
  assign _T_97407 = _T_90415 ? _T_97405 : 16'h0; // @[Mux.scala 19:72:@41687.4]
  assign _T_97408 = _T_97152 | _T_97169; // @[Mux.scala 19:72:@41688.4]
  assign _T_97409 = _T_97408 | _T_97186; // @[Mux.scala 19:72:@41689.4]
  assign _T_97410 = _T_97409 | _T_97203; // @[Mux.scala 19:72:@41690.4]
  assign _T_97411 = _T_97410 | _T_97220; // @[Mux.scala 19:72:@41691.4]
  assign _T_97412 = _T_97411 | _T_97237; // @[Mux.scala 19:72:@41692.4]
  assign _T_97413 = _T_97412 | _T_97254; // @[Mux.scala 19:72:@41693.4]
  assign _T_97414 = _T_97413 | _T_97271; // @[Mux.scala 19:72:@41694.4]
  assign _T_97415 = _T_97414 | _T_97288; // @[Mux.scala 19:72:@41695.4]
  assign _T_97416 = _T_97415 | _T_97305; // @[Mux.scala 19:72:@41696.4]
  assign _T_97417 = _T_97416 | _T_97322; // @[Mux.scala 19:72:@41697.4]
  assign _T_97418 = _T_97417 | _T_97339; // @[Mux.scala 19:72:@41698.4]
  assign _T_97419 = _T_97418 | _T_97356; // @[Mux.scala 19:72:@41699.4]
  assign _T_97420 = _T_97419 | _T_97373; // @[Mux.scala 19:72:@41700.4]
  assign _T_97421 = _T_97420 | _T_97390; // @[Mux.scala 19:72:@41701.4]
  assign _T_97422 = _T_97421 | _T_97407; // @[Mux.scala 19:72:@41702.4]
  assign outputPriorityPorts_0_0 = _T_97422[0]; // @[Mux.scala 19:72:@41706.4]
  assign outputPriorityPorts_0_1 = _T_97422[1]; // @[Mux.scala 19:72:@41708.4]
  assign outputPriorityPorts_0_2 = _T_97422[2]; // @[Mux.scala 19:72:@41710.4]
  assign outputPriorityPorts_0_3 = _T_97422[3]; // @[Mux.scala 19:72:@41712.4]
  assign outputPriorityPorts_0_4 = _T_97422[4]; // @[Mux.scala 19:72:@41714.4]
  assign outputPriorityPorts_0_5 = _T_97422[5]; // @[Mux.scala 19:72:@41716.4]
  assign outputPriorityPorts_0_6 = _T_97422[6]; // @[Mux.scala 19:72:@41718.4]
  assign outputPriorityPorts_0_7 = _T_97422[7]; // @[Mux.scala 19:72:@41720.4]
  assign outputPriorityPorts_0_8 = _T_97422[8]; // @[Mux.scala 19:72:@41722.4]
  assign outputPriorityPorts_0_9 = _T_97422[9]; // @[Mux.scala 19:72:@41724.4]
  assign outputPriorityPorts_0_10 = _T_97422[10]; // @[Mux.scala 19:72:@41726.4]
  assign outputPriorityPorts_0_11 = _T_97422[11]; // @[Mux.scala 19:72:@41728.4]
  assign outputPriorityPorts_0_12 = _T_97422[12]; // @[Mux.scala 19:72:@41730.4]
  assign outputPriorityPorts_0_13 = _T_97422[13]; // @[Mux.scala 19:72:@41732.4]
  assign outputPriorityPorts_0_14 = _T_97422[14]; // @[Mux.scala 19:72:@41734.4]
  assign outputPriorityPorts_0_15 = _T_97422[15]; // @[Mux.scala 19:72:@41736.4]
  assign _T_97565 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41758.6]
  assign _GEN_2114 = _T_97565 ? io_addrFromLoadPorts_0 : addrQ_0; // @[LoadQueue.scala 314:36:@41762.6]
  assign _GEN_2115 = _T_97565 ? 1'h1 : addrKnown_0; // @[LoadQueue.scala 314:36:@41762.6]
  assign _GEN_2116 = initBits_0 ? 1'h0 : _GEN_2115; // @[LoadQueue.scala 308:34:@41754.4]
  assign _GEN_2117 = initBits_0 ? addrQ_0 : _GEN_2114; // @[LoadQueue.scala 308:34:@41754.4]
  assign _T_97580 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41771.6]
  assign _GEN_2118 = _T_97580 ? io_addrFromLoadPorts_0 : addrQ_1; // @[LoadQueue.scala 314:36:@41775.6]
  assign _GEN_2119 = _T_97580 ? 1'h1 : addrKnown_1; // @[LoadQueue.scala 314:36:@41775.6]
  assign _GEN_2120 = initBits_1 ? 1'h0 : _GEN_2119; // @[LoadQueue.scala 308:34:@41767.4]
  assign _GEN_2121 = initBits_1 ? addrQ_1 : _GEN_2118; // @[LoadQueue.scala 308:34:@41767.4]
  assign _T_97595 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41784.6]
  assign _GEN_2122 = _T_97595 ? io_addrFromLoadPorts_0 : addrQ_2; // @[LoadQueue.scala 314:36:@41788.6]
  assign _GEN_2123 = _T_97595 ? 1'h1 : addrKnown_2; // @[LoadQueue.scala 314:36:@41788.6]
  assign _GEN_2124 = initBits_2 ? 1'h0 : _GEN_2123; // @[LoadQueue.scala 308:34:@41780.4]
  assign _GEN_2125 = initBits_2 ? addrQ_2 : _GEN_2122; // @[LoadQueue.scala 308:34:@41780.4]
  assign _T_97610 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41797.6]
  assign _GEN_2126 = _T_97610 ? io_addrFromLoadPorts_0 : addrQ_3; // @[LoadQueue.scala 314:36:@41801.6]
  assign _GEN_2127 = _T_97610 ? 1'h1 : addrKnown_3; // @[LoadQueue.scala 314:36:@41801.6]
  assign _GEN_2128 = initBits_3 ? 1'h0 : _GEN_2127; // @[LoadQueue.scala 308:34:@41793.4]
  assign _GEN_2129 = initBits_3 ? addrQ_3 : _GEN_2126; // @[LoadQueue.scala 308:34:@41793.4]
  assign _T_97625 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41810.6]
  assign _GEN_2130 = _T_97625 ? io_addrFromLoadPorts_0 : addrQ_4; // @[LoadQueue.scala 314:36:@41814.6]
  assign _GEN_2131 = _T_97625 ? 1'h1 : addrKnown_4; // @[LoadQueue.scala 314:36:@41814.6]
  assign _GEN_2132 = initBits_4 ? 1'h0 : _GEN_2131; // @[LoadQueue.scala 308:34:@41806.4]
  assign _GEN_2133 = initBits_4 ? addrQ_4 : _GEN_2130; // @[LoadQueue.scala 308:34:@41806.4]
  assign _T_97640 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41823.6]
  assign _GEN_2134 = _T_97640 ? io_addrFromLoadPorts_0 : addrQ_5; // @[LoadQueue.scala 314:36:@41827.6]
  assign _GEN_2135 = _T_97640 ? 1'h1 : addrKnown_5; // @[LoadQueue.scala 314:36:@41827.6]
  assign _GEN_2136 = initBits_5 ? 1'h0 : _GEN_2135; // @[LoadQueue.scala 308:34:@41819.4]
  assign _GEN_2137 = initBits_5 ? addrQ_5 : _GEN_2134; // @[LoadQueue.scala 308:34:@41819.4]
  assign _T_97655 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41836.6]
  assign _GEN_2138 = _T_97655 ? io_addrFromLoadPorts_0 : addrQ_6; // @[LoadQueue.scala 314:36:@41840.6]
  assign _GEN_2139 = _T_97655 ? 1'h1 : addrKnown_6; // @[LoadQueue.scala 314:36:@41840.6]
  assign _GEN_2140 = initBits_6 ? 1'h0 : _GEN_2139; // @[LoadQueue.scala 308:34:@41832.4]
  assign _GEN_2141 = initBits_6 ? addrQ_6 : _GEN_2138; // @[LoadQueue.scala 308:34:@41832.4]
  assign _T_97670 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41849.6]
  assign _GEN_2142 = _T_97670 ? io_addrFromLoadPorts_0 : addrQ_7; // @[LoadQueue.scala 314:36:@41853.6]
  assign _GEN_2143 = _T_97670 ? 1'h1 : addrKnown_7; // @[LoadQueue.scala 314:36:@41853.6]
  assign _GEN_2144 = initBits_7 ? 1'h0 : _GEN_2143; // @[LoadQueue.scala 308:34:@41845.4]
  assign _GEN_2145 = initBits_7 ? addrQ_7 : _GEN_2142; // @[LoadQueue.scala 308:34:@41845.4]
  assign _T_97685 = inputPriorityPorts_0_8 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41862.6]
  assign _GEN_2146 = _T_97685 ? io_addrFromLoadPorts_0 : addrQ_8; // @[LoadQueue.scala 314:36:@41866.6]
  assign _GEN_2147 = _T_97685 ? 1'h1 : addrKnown_8; // @[LoadQueue.scala 314:36:@41866.6]
  assign _GEN_2148 = initBits_8 ? 1'h0 : _GEN_2147; // @[LoadQueue.scala 308:34:@41858.4]
  assign _GEN_2149 = initBits_8 ? addrQ_8 : _GEN_2146; // @[LoadQueue.scala 308:34:@41858.4]
  assign _T_97700 = inputPriorityPorts_0_9 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41875.6]
  assign _GEN_2150 = _T_97700 ? io_addrFromLoadPorts_0 : addrQ_9; // @[LoadQueue.scala 314:36:@41879.6]
  assign _GEN_2151 = _T_97700 ? 1'h1 : addrKnown_9; // @[LoadQueue.scala 314:36:@41879.6]
  assign _GEN_2152 = initBits_9 ? 1'h0 : _GEN_2151; // @[LoadQueue.scala 308:34:@41871.4]
  assign _GEN_2153 = initBits_9 ? addrQ_9 : _GEN_2150; // @[LoadQueue.scala 308:34:@41871.4]
  assign _T_97715 = inputPriorityPorts_0_10 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41888.6]
  assign _GEN_2154 = _T_97715 ? io_addrFromLoadPorts_0 : addrQ_10; // @[LoadQueue.scala 314:36:@41892.6]
  assign _GEN_2155 = _T_97715 ? 1'h1 : addrKnown_10; // @[LoadQueue.scala 314:36:@41892.6]
  assign _GEN_2156 = initBits_10 ? 1'h0 : _GEN_2155; // @[LoadQueue.scala 308:34:@41884.4]
  assign _GEN_2157 = initBits_10 ? addrQ_10 : _GEN_2154; // @[LoadQueue.scala 308:34:@41884.4]
  assign _T_97730 = inputPriorityPorts_0_11 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41901.6]
  assign _GEN_2158 = _T_97730 ? io_addrFromLoadPorts_0 : addrQ_11; // @[LoadQueue.scala 314:36:@41905.6]
  assign _GEN_2159 = _T_97730 ? 1'h1 : addrKnown_11; // @[LoadQueue.scala 314:36:@41905.6]
  assign _GEN_2160 = initBits_11 ? 1'h0 : _GEN_2159; // @[LoadQueue.scala 308:34:@41897.4]
  assign _GEN_2161 = initBits_11 ? addrQ_11 : _GEN_2158; // @[LoadQueue.scala 308:34:@41897.4]
  assign _T_97745 = inputPriorityPorts_0_12 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41914.6]
  assign _GEN_2162 = _T_97745 ? io_addrFromLoadPorts_0 : addrQ_12; // @[LoadQueue.scala 314:36:@41918.6]
  assign _GEN_2163 = _T_97745 ? 1'h1 : addrKnown_12; // @[LoadQueue.scala 314:36:@41918.6]
  assign _GEN_2164 = initBits_12 ? 1'h0 : _GEN_2163; // @[LoadQueue.scala 308:34:@41910.4]
  assign _GEN_2165 = initBits_12 ? addrQ_12 : _GEN_2162; // @[LoadQueue.scala 308:34:@41910.4]
  assign _T_97760 = inputPriorityPorts_0_13 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41927.6]
  assign _GEN_2166 = _T_97760 ? io_addrFromLoadPorts_0 : addrQ_13; // @[LoadQueue.scala 314:36:@41931.6]
  assign _GEN_2167 = _T_97760 ? 1'h1 : addrKnown_13; // @[LoadQueue.scala 314:36:@41931.6]
  assign _GEN_2168 = initBits_13 ? 1'h0 : _GEN_2167; // @[LoadQueue.scala 308:34:@41923.4]
  assign _GEN_2169 = initBits_13 ? addrQ_13 : _GEN_2166; // @[LoadQueue.scala 308:34:@41923.4]
  assign _T_97775 = inputPriorityPorts_0_14 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41940.6]
  assign _GEN_2170 = _T_97775 ? io_addrFromLoadPorts_0 : addrQ_14; // @[LoadQueue.scala 314:36:@41944.6]
  assign _GEN_2171 = _T_97775 ? 1'h1 : addrKnown_14; // @[LoadQueue.scala 314:36:@41944.6]
  assign _GEN_2172 = initBits_14 ? 1'h0 : _GEN_2171; // @[LoadQueue.scala 308:34:@41936.4]
  assign _GEN_2173 = initBits_14 ? addrQ_14 : _GEN_2170; // @[LoadQueue.scala 308:34:@41936.4]
  assign _T_97790 = inputPriorityPorts_0_15 & io_loadAddrEnable_0; // @[LoadQueue.scala 313:47:@41953.6]
  assign _GEN_2174 = _T_97790 ? io_addrFromLoadPorts_0 : addrQ_15; // @[LoadQueue.scala 314:36:@41957.6]
  assign _GEN_2175 = _T_97790 ? 1'h1 : addrKnown_15; // @[LoadQueue.scala 314:36:@41957.6]
  assign _GEN_2176 = initBits_15 ? 1'h0 : _GEN_2175; // @[LoadQueue.scala 308:34:@41949.4]
  assign _GEN_2177 = initBits_15 ? addrQ_15 : _GEN_2174; // @[LoadQueue.scala 308:34:@41949.4]
  assign _T_97825 = outputPriorityPorts_0_0 & dataKnown_0; // @[LoadQueue.scala 326:108:@41963.4]
  assign _T_97827 = loadCompleted_0 == 1'h0; // @[LoadQueue.scala 327:34:@41964.4]
  assign _T_97828 = _T_97825 & _T_97827; // @[LoadQueue.scala 327:31:@41965.4]
  assign loadCompleting_0 = _T_97828 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@41966.4]
  assign _T_97839 = outputPriorityPorts_0_1 & dataKnown_1; // @[LoadQueue.scala 326:108:@41971.4]
  assign _T_97841 = loadCompleted_1 == 1'h0; // @[LoadQueue.scala 327:34:@41972.4]
  assign _T_97842 = _T_97839 & _T_97841; // @[LoadQueue.scala 327:31:@41973.4]
  assign loadCompleting_1 = _T_97842 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@41974.4]
  assign _T_97853 = outputPriorityPorts_0_2 & dataKnown_2; // @[LoadQueue.scala 326:108:@41979.4]
  assign _T_97855 = loadCompleted_2 == 1'h0; // @[LoadQueue.scala 327:34:@41980.4]
  assign _T_97856 = _T_97853 & _T_97855; // @[LoadQueue.scala 327:31:@41981.4]
  assign loadCompleting_2 = _T_97856 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@41982.4]
  assign _T_97867 = outputPriorityPorts_0_3 & dataKnown_3; // @[LoadQueue.scala 326:108:@41987.4]
  assign _T_97869 = loadCompleted_3 == 1'h0; // @[LoadQueue.scala 327:34:@41988.4]
  assign _T_97870 = _T_97867 & _T_97869; // @[LoadQueue.scala 327:31:@41989.4]
  assign loadCompleting_3 = _T_97870 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@41990.4]
  assign _T_97881 = outputPriorityPorts_0_4 & dataKnown_4; // @[LoadQueue.scala 326:108:@41995.4]
  assign _T_97883 = loadCompleted_4 == 1'h0; // @[LoadQueue.scala 327:34:@41996.4]
  assign _T_97884 = _T_97881 & _T_97883; // @[LoadQueue.scala 327:31:@41997.4]
  assign loadCompleting_4 = _T_97884 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@41998.4]
  assign _T_97895 = outputPriorityPorts_0_5 & dataKnown_5; // @[LoadQueue.scala 326:108:@42003.4]
  assign _T_97897 = loadCompleted_5 == 1'h0; // @[LoadQueue.scala 327:34:@42004.4]
  assign _T_97898 = _T_97895 & _T_97897; // @[LoadQueue.scala 327:31:@42005.4]
  assign loadCompleting_5 = _T_97898 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42006.4]
  assign _T_97909 = outputPriorityPorts_0_6 & dataKnown_6; // @[LoadQueue.scala 326:108:@42011.4]
  assign _T_97911 = loadCompleted_6 == 1'h0; // @[LoadQueue.scala 327:34:@42012.4]
  assign _T_97912 = _T_97909 & _T_97911; // @[LoadQueue.scala 327:31:@42013.4]
  assign loadCompleting_6 = _T_97912 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42014.4]
  assign _T_97923 = outputPriorityPorts_0_7 & dataKnown_7; // @[LoadQueue.scala 326:108:@42019.4]
  assign _T_97925 = loadCompleted_7 == 1'h0; // @[LoadQueue.scala 327:34:@42020.4]
  assign _T_97926 = _T_97923 & _T_97925; // @[LoadQueue.scala 327:31:@42021.4]
  assign loadCompleting_7 = _T_97926 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42022.4]
  assign _T_97937 = outputPriorityPorts_0_8 & dataKnown_8; // @[LoadQueue.scala 326:108:@42027.4]
  assign _T_97939 = loadCompleted_8 == 1'h0; // @[LoadQueue.scala 327:34:@42028.4]
  assign _T_97940 = _T_97937 & _T_97939; // @[LoadQueue.scala 327:31:@42029.4]
  assign loadCompleting_8 = _T_97940 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42030.4]
  assign _T_97951 = outputPriorityPorts_0_9 & dataKnown_9; // @[LoadQueue.scala 326:108:@42035.4]
  assign _T_97953 = loadCompleted_9 == 1'h0; // @[LoadQueue.scala 327:34:@42036.4]
  assign _T_97954 = _T_97951 & _T_97953; // @[LoadQueue.scala 327:31:@42037.4]
  assign loadCompleting_9 = _T_97954 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42038.4]
  assign _T_97965 = outputPriorityPorts_0_10 & dataKnown_10; // @[LoadQueue.scala 326:108:@42043.4]
  assign _T_97967 = loadCompleted_10 == 1'h0; // @[LoadQueue.scala 327:34:@42044.4]
  assign _T_97968 = _T_97965 & _T_97967; // @[LoadQueue.scala 327:31:@42045.4]
  assign loadCompleting_10 = _T_97968 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42046.4]
  assign _T_97979 = outputPriorityPorts_0_11 & dataKnown_11; // @[LoadQueue.scala 326:108:@42051.4]
  assign _T_97981 = loadCompleted_11 == 1'h0; // @[LoadQueue.scala 327:34:@42052.4]
  assign _T_97982 = _T_97979 & _T_97981; // @[LoadQueue.scala 327:31:@42053.4]
  assign loadCompleting_11 = _T_97982 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42054.4]
  assign _T_97993 = outputPriorityPorts_0_12 & dataKnown_12; // @[LoadQueue.scala 326:108:@42059.4]
  assign _T_97995 = loadCompleted_12 == 1'h0; // @[LoadQueue.scala 327:34:@42060.4]
  assign _T_97996 = _T_97993 & _T_97995; // @[LoadQueue.scala 327:31:@42061.4]
  assign loadCompleting_12 = _T_97996 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42062.4]
  assign _T_98007 = outputPriorityPorts_0_13 & dataKnown_13; // @[LoadQueue.scala 326:108:@42067.4]
  assign _T_98009 = loadCompleted_13 == 1'h0; // @[LoadQueue.scala 327:34:@42068.4]
  assign _T_98010 = _T_98007 & _T_98009; // @[LoadQueue.scala 327:31:@42069.4]
  assign loadCompleting_13 = _T_98010 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42070.4]
  assign _T_98021 = outputPriorityPorts_0_14 & dataKnown_14; // @[LoadQueue.scala 326:108:@42075.4]
  assign _T_98023 = loadCompleted_14 == 1'h0; // @[LoadQueue.scala 327:34:@42076.4]
  assign _T_98024 = _T_98021 & _T_98023; // @[LoadQueue.scala 327:31:@42077.4]
  assign loadCompleting_14 = _T_98024 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42078.4]
  assign _T_98035 = outputPriorityPorts_0_15 & dataKnown_15; // @[LoadQueue.scala 326:108:@42083.4]
  assign _T_98037 = loadCompleted_15 == 1'h0; // @[LoadQueue.scala 327:34:@42084.4]
  assign _T_98038 = _T_98035 & _T_98037; // @[LoadQueue.scala 327:31:@42085.4]
  assign loadCompleting_15 = _T_98038 & io_loadPorts_0_ready; // @[LoadQueue.scala 327:63:@42086.4]
  assign _GEN_2178 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[LoadQueue.scala 337:46:@42095.6]
  assign _GEN_2179 = initBits_0 ? 1'h0 : _GEN_2178; // @[LoadQueue.scala 335:34:@42091.4]
  assign _GEN_2180 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[LoadQueue.scala 337:46:@42102.6]
  assign _GEN_2181 = initBits_1 ? 1'h0 : _GEN_2180; // @[LoadQueue.scala 335:34:@42098.4]
  assign _GEN_2182 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[LoadQueue.scala 337:46:@42109.6]
  assign _GEN_2183 = initBits_2 ? 1'h0 : _GEN_2182; // @[LoadQueue.scala 335:34:@42105.4]
  assign _GEN_2184 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[LoadQueue.scala 337:46:@42116.6]
  assign _GEN_2185 = initBits_3 ? 1'h0 : _GEN_2184; // @[LoadQueue.scala 335:34:@42112.4]
  assign _GEN_2186 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[LoadQueue.scala 337:46:@42123.6]
  assign _GEN_2187 = initBits_4 ? 1'h0 : _GEN_2186; // @[LoadQueue.scala 335:34:@42119.4]
  assign _GEN_2188 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[LoadQueue.scala 337:46:@42130.6]
  assign _GEN_2189 = initBits_5 ? 1'h0 : _GEN_2188; // @[LoadQueue.scala 335:34:@42126.4]
  assign _GEN_2190 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[LoadQueue.scala 337:46:@42137.6]
  assign _GEN_2191 = initBits_6 ? 1'h0 : _GEN_2190; // @[LoadQueue.scala 335:34:@42133.4]
  assign _GEN_2192 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[LoadQueue.scala 337:46:@42144.6]
  assign _GEN_2193 = initBits_7 ? 1'h0 : _GEN_2192; // @[LoadQueue.scala 335:34:@42140.4]
  assign _GEN_2194 = loadCompleting_8 ? 1'h1 : loadCompleted_8; // @[LoadQueue.scala 337:46:@42151.6]
  assign _GEN_2195 = initBits_8 ? 1'h0 : _GEN_2194; // @[LoadQueue.scala 335:34:@42147.4]
  assign _GEN_2196 = loadCompleting_9 ? 1'h1 : loadCompleted_9; // @[LoadQueue.scala 337:46:@42158.6]
  assign _GEN_2197 = initBits_9 ? 1'h0 : _GEN_2196; // @[LoadQueue.scala 335:34:@42154.4]
  assign _GEN_2198 = loadCompleting_10 ? 1'h1 : loadCompleted_10; // @[LoadQueue.scala 337:46:@42165.6]
  assign _GEN_2199 = initBits_10 ? 1'h0 : _GEN_2198; // @[LoadQueue.scala 335:34:@42161.4]
  assign _GEN_2200 = loadCompleting_11 ? 1'h1 : loadCompleted_11; // @[LoadQueue.scala 337:46:@42172.6]
  assign _GEN_2201 = initBits_11 ? 1'h0 : _GEN_2200; // @[LoadQueue.scala 335:34:@42168.4]
  assign _GEN_2202 = loadCompleting_12 ? 1'h1 : loadCompleted_12; // @[LoadQueue.scala 337:46:@42179.6]
  assign _GEN_2203 = initBits_12 ? 1'h0 : _GEN_2202; // @[LoadQueue.scala 335:34:@42175.4]
  assign _GEN_2204 = loadCompleting_13 ? 1'h1 : loadCompleted_13; // @[LoadQueue.scala 337:46:@42186.6]
  assign _GEN_2205 = initBits_13 ? 1'h0 : _GEN_2204; // @[LoadQueue.scala 335:34:@42182.4]
  assign _GEN_2206 = loadCompleting_14 ? 1'h1 : loadCompleted_14; // @[LoadQueue.scala 337:46:@42193.6]
  assign _GEN_2207 = initBits_14 ? 1'h0 : _GEN_2206; // @[LoadQueue.scala 335:34:@42189.4]
  assign _GEN_2208 = loadCompleting_15 ? 1'h1 : loadCompleted_15; // @[LoadQueue.scala 337:46:@42200.6]
  assign _GEN_2209 = initBits_15 ? 1'h0 : _GEN_2208; // @[LoadQueue.scala 335:34:@42196.4]
  assign _T_98169 = _T_97828 | _T_97842; // @[LoadQueue.scala 348:24:@42269.4]
  assign _T_98170 = _T_98169 | _T_97856; // @[LoadQueue.scala 348:24:@42270.4]
  assign _T_98171 = _T_98170 | _T_97870; // @[LoadQueue.scala 348:24:@42271.4]
  assign _T_98172 = _T_98171 | _T_97884; // @[LoadQueue.scala 348:24:@42272.4]
  assign _T_98173 = _T_98172 | _T_97898; // @[LoadQueue.scala 348:24:@42273.4]
  assign _T_98174 = _T_98173 | _T_97912; // @[LoadQueue.scala 348:24:@42274.4]
  assign _T_98175 = _T_98174 | _T_97926; // @[LoadQueue.scala 348:24:@42275.4]
  assign _T_98176 = _T_98175 | _T_97940; // @[LoadQueue.scala 348:24:@42276.4]
  assign _T_98177 = _T_98176 | _T_97954; // @[LoadQueue.scala 348:24:@42277.4]
  assign _T_98178 = _T_98177 | _T_97968; // @[LoadQueue.scala 348:24:@42278.4]
  assign _T_98179 = _T_98178 | _T_97982; // @[LoadQueue.scala 348:24:@42279.4]
  assign _T_98180 = _T_98179 | _T_97996; // @[LoadQueue.scala 348:24:@42280.4]
  assign _T_98181 = _T_98180 | _T_98010; // @[LoadQueue.scala 348:24:@42281.4]
  assign _T_98182 = _T_98181 | _T_98024; // @[LoadQueue.scala 348:24:@42282.4]
  assign _T_98183 = _T_98182 | _T_98038; // @[LoadQueue.scala 348:24:@42283.4]
  assign _T_98200 = _T_98024 ? 4'he : 4'hf; // @[Mux.scala 31:69:@42285.6]
  assign _T_98201 = _T_98010 ? 4'hd : _T_98200; // @[Mux.scala 31:69:@42286.6]
  assign _T_98202 = _T_97996 ? 4'hc : _T_98201; // @[Mux.scala 31:69:@42287.6]
  assign _T_98203 = _T_97982 ? 4'hb : _T_98202; // @[Mux.scala 31:69:@42288.6]
  assign _T_98204 = _T_97968 ? 4'ha : _T_98203; // @[Mux.scala 31:69:@42289.6]
  assign _T_98205 = _T_97954 ? 4'h9 : _T_98204; // @[Mux.scala 31:69:@42290.6]
  assign _T_98206 = _T_97940 ? 4'h8 : _T_98205; // @[Mux.scala 31:69:@42291.6]
  assign _T_98207 = _T_97926 ? 4'h7 : _T_98206; // @[Mux.scala 31:69:@42292.6]
  assign _T_98208 = _T_97912 ? 4'h6 : _T_98207; // @[Mux.scala 31:69:@42293.6]
  assign _T_98209 = _T_97898 ? 4'h5 : _T_98208; // @[Mux.scala 31:69:@42294.6]
  assign _T_98210 = _T_97884 ? 4'h4 : _T_98209; // @[Mux.scala 31:69:@42295.6]
  assign _T_98211 = _T_97870 ? 4'h3 : _T_98210; // @[Mux.scala 31:69:@42296.6]
  assign _T_98212 = _T_97856 ? 4'h2 : _T_98211; // @[Mux.scala 31:69:@42297.6]
  assign _T_98213 = _T_97842 ? 4'h1 : _T_98212; // @[Mux.scala 31:69:@42298.6]
  assign _T_98214 = _T_97828 ? 4'h0 : _T_98213; // @[Mux.scala 31:69:@42299.6]
  assign _GEN_2211 = 4'h1 == _T_98214 ? dataQ_1 : dataQ_0; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2212 = 4'h2 == _T_98214 ? dataQ_2 : _GEN_2211; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2213 = 4'h3 == _T_98214 ? dataQ_3 : _GEN_2212; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2214 = 4'h4 == _T_98214 ? dataQ_4 : _GEN_2213; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2215 = 4'h5 == _T_98214 ? dataQ_5 : _GEN_2214; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2216 = 4'h6 == _T_98214 ? dataQ_6 : _GEN_2215; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2217 = 4'h7 == _T_98214 ? dataQ_7 : _GEN_2216; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2218 = 4'h8 == _T_98214 ? dataQ_8 : _GEN_2217; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2219 = 4'h9 == _T_98214 ? dataQ_9 : _GEN_2218; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2220 = 4'ha == _T_98214 ? dataQ_10 : _GEN_2219; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2221 = 4'hb == _T_98214 ? dataQ_11 : _GEN_2220; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2222 = 4'hc == _T_98214 ? dataQ_12 : _GEN_2221; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2223 = 4'hd == _T_98214 ? dataQ_13 : _GEN_2222; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2224 = 4'he == _T_98214 ? dataQ_14 : _GEN_2223; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2225 = 4'hf == _T_98214 ? dataQ_15 : _GEN_2224; // @[LoadQueue.scala 349:37:@42300.6]
  assign _GEN_2229 = 4'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2230 = 4'h2 == head ? loadCompleted_2 : _GEN_2229; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2231 = 4'h3 == head ? loadCompleted_3 : _GEN_2230; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2232 = 4'h4 == head ? loadCompleted_4 : _GEN_2231; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2233 = 4'h5 == head ? loadCompleted_5 : _GEN_2232; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2234 = 4'h6 == head ? loadCompleted_6 : _GEN_2233; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2235 = 4'h7 == head ? loadCompleted_7 : _GEN_2234; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2236 = 4'h8 == head ? loadCompleted_8 : _GEN_2235; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2237 = 4'h9 == head ? loadCompleted_9 : _GEN_2236; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2238 = 4'ha == head ? loadCompleted_10 : _GEN_2237; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2239 = 4'hb == head ? loadCompleted_11 : _GEN_2238; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2240 = 4'hc == head ? loadCompleted_12 : _GEN_2239; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2241 = 4'hd == head ? loadCompleted_13 : _GEN_2240; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2242 = 4'he == head ? loadCompleted_14 : _GEN_2241; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2243 = 4'hf == head ? loadCompleted_15 : _GEN_2242; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2245 = 4'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2246 = 4'h2 == head ? loadCompleting_2 : _GEN_2245; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2247 = 4'h3 == head ? loadCompleting_3 : _GEN_2246; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2248 = 4'h4 == head ? loadCompleting_4 : _GEN_2247; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2249 = 4'h5 == head ? loadCompleting_5 : _GEN_2248; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2250 = 4'h6 == head ? loadCompleting_6 : _GEN_2249; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2251 = 4'h7 == head ? loadCompleting_7 : _GEN_2250; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2252 = 4'h8 == head ? loadCompleting_8 : _GEN_2251; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2253 = 4'h9 == head ? loadCompleting_9 : _GEN_2252; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2254 = 4'ha == head ? loadCompleting_10 : _GEN_2253; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2255 = 4'hb == head ? loadCompleting_11 : _GEN_2254; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2256 = 4'hc == head ? loadCompleting_12 : _GEN_2255; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2257 = 4'hd == head ? loadCompleting_13 : _GEN_2256; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2258 = 4'he == head ? loadCompleting_14 : _GEN_2257; // @[LoadQueue.scala 363:29:@42307.4]
  assign _GEN_2259 = 4'hf == head ? loadCompleting_15 : _GEN_2258; // @[LoadQueue.scala 363:29:@42307.4]
  assign _T_98225 = _GEN_2243 | _GEN_2259; // @[LoadQueue.scala 363:29:@42307.4]
  assign _T_98226 = head != tail; // @[LoadQueue.scala 363:63:@42308.4]
  assign _T_98228 = io_loadEmpty == 1'h0; // @[LoadQueue.scala 363:75:@42309.4]
  assign _T_98229 = _T_98226 | _T_98228; // @[LoadQueue.scala 363:72:@42310.4]
  assign _T_98230 = _T_98225 & _T_98229; // @[LoadQueue.scala 363:54:@42311.4]
  assign _T_98233 = head + 4'h1; // @[util.scala 10:8:@42313.6]
  assign _GEN_64 = _T_98233 % 5'h10; // @[util.scala 10:14:@42314.6]
  assign _T_98234 = _GEN_64[4:0]; // @[util.scala 10:14:@42314.6]
  assign _GEN_2260 = _T_98230 ? _T_98234 : {{1'd0}, head}; // @[LoadQueue.scala 363:91:@42312.4]
  assign _GEN_2358 = {{3'd0}, io_bbNumLoads}; // @[util.scala 10:8:@42318.6]
  assign _T_98236 = tail + _GEN_2358; // @[util.scala 10:8:@42318.6]
  assign _GEN_65 = _T_98236 % 5'h10; // @[util.scala 10:14:@42319.6]
  assign _T_98237 = _GEN_65[4:0]; // @[util.scala 10:14:@42319.6]
  assign _GEN_2261 = io_bbStart ? _T_98237 : {{1'd0}, tail}; // @[LoadQueue.scala 367:20:@42317.4]
  assign _T_98239 = allocatedEntries_0 == 1'h0; // @[LoadQueue.scala 371:82:@42322.4]
  assign _T_98240 = loadCompleted_0 | _T_98239; // @[LoadQueue.scala 371:79:@42323.4]
  assign _T_98242 = allocatedEntries_1 == 1'h0; // @[LoadQueue.scala 371:82:@42324.4]
  assign _T_98243 = loadCompleted_1 | _T_98242; // @[LoadQueue.scala 371:79:@42325.4]
  assign _T_98245 = allocatedEntries_2 == 1'h0; // @[LoadQueue.scala 371:82:@42326.4]
  assign _T_98246 = loadCompleted_2 | _T_98245; // @[LoadQueue.scala 371:79:@42327.4]
  assign _T_98248 = allocatedEntries_3 == 1'h0; // @[LoadQueue.scala 371:82:@42328.4]
  assign _T_98249 = loadCompleted_3 | _T_98248; // @[LoadQueue.scala 371:79:@42329.4]
  assign _T_98251 = allocatedEntries_4 == 1'h0; // @[LoadQueue.scala 371:82:@42330.4]
  assign _T_98252 = loadCompleted_4 | _T_98251; // @[LoadQueue.scala 371:79:@42331.4]
  assign _T_98254 = allocatedEntries_5 == 1'h0; // @[LoadQueue.scala 371:82:@42332.4]
  assign _T_98255 = loadCompleted_5 | _T_98254; // @[LoadQueue.scala 371:79:@42333.4]
  assign _T_98257 = allocatedEntries_6 == 1'h0; // @[LoadQueue.scala 371:82:@42334.4]
  assign _T_98258 = loadCompleted_6 | _T_98257; // @[LoadQueue.scala 371:79:@42335.4]
  assign _T_98260 = allocatedEntries_7 == 1'h0; // @[LoadQueue.scala 371:82:@42336.4]
  assign _T_98261 = loadCompleted_7 | _T_98260; // @[LoadQueue.scala 371:79:@42337.4]
  assign _T_98263 = allocatedEntries_8 == 1'h0; // @[LoadQueue.scala 371:82:@42338.4]
  assign _T_98264 = loadCompleted_8 | _T_98263; // @[LoadQueue.scala 371:79:@42339.4]
  assign _T_98266 = allocatedEntries_9 == 1'h0; // @[LoadQueue.scala 371:82:@42340.4]
  assign _T_98267 = loadCompleted_9 | _T_98266; // @[LoadQueue.scala 371:79:@42341.4]
  assign _T_98269 = allocatedEntries_10 == 1'h0; // @[LoadQueue.scala 371:82:@42342.4]
  assign _T_98270 = loadCompleted_10 | _T_98269; // @[LoadQueue.scala 371:79:@42343.4]
  assign _T_98272 = allocatedEntries_11 == 1'h0; // @[LoadQueue.scala 371:82:@42344.4]
  assign _T_98273 = loadCompleted_11 | _T_98272; // @[LoadQueue.scala 371:79:@42345.4]
  assign _T_98275 = allocatedEntries_12 == 1'h0; // @[LoadQueue.scala 371:82:@42346.4]
  assign _T_98276 = loadCompleted_12 | _T_98275; // @[LoadQueue.scala 371:79:@42347.4]
  assign _T_98278 = allocatedEntries_13 == 1'h0; // @[LoadQueue.scala 371:82:@42348.4]
  assign _T_98279 = loadCompleted_13 | _T_98278; // @[LoadQueue.scala 371:79:@42349.4]
  assign _T_98281 = allocatedEntries_14 == 1'h0; // @[LoadQueue.scala 371:82:@42350.4]
  assign _T_98282 = loadCompleted_14 | _T_98281; // @[LoadQueue.scala 371:79:@42351.4]
  assign _T_98284 = allocatedEntries_15 == 1'h0; // @[LoadQueue.scala 371:82:@42352.4]
  assign _T_98285 = loadCompleted_15 | _T_98284; // @[LoadQueue.scala 371:79:@42353.4]
  assign _T_98310 = _T_98240 & _T_98243; // @[LoadQueue.scala 371:96:@42372.4]
  assign _T_98311 = _T_98310 & _T_98246; // @[LoadQueue.scala 371:96:@42373.4]
  assign _T_98312 = _T_98311 & _T_98249; // @[LoadQueue.scala 371:96:@42374.4]
  assign _T_98313 = _T_98312 & _T_98252; // @[LoadQueue.scala 371:96:@42375.4]
  assign _T_98314 = _T_98313 & _T_98255; // @[LoadQueue.scala 371:96:@42376.4]
  assign _T_98315 = _T_98314 & _T_98258; // @[LoadQueue.scala 371:96:@42377.4]
  assign _T_98316 = _T_98315 & _T_98261; // @[LoadQueue.scala 371:96:@42378.4]
  assign _T_98317 = _T_98316 & _T_98264; // @[LoadQueue.scala 371:96:@42379.4]
  assign _T_98318 = _T_98317 & _T_98267; // @[LoadQueue.scala 371:96:@42380.4]
  assign _T_98319 = _T_98318 & _T_98270; // @[LoadQueue.scala 371:96:@42381.4]
  assign _T_98320 = _T_98319 & _T_98273; // @[LoadQueue.scala 371:96:@42382.4]
  assign _T_98321 = _T_98320 & _T_98276; // @[LoadQueue.scala 371:96:@42383.4]
  assign _T_98322 = _T_98321 & _T_98279; // @[LoadQueue.scala 371:96:@42384.4]
  assign _T_98323 = _T_98322 & _T_98282; // @[LoadQueue.scala 371:96:@42385.4]
  assign io_loadTail = tail; // @[LoadQueue.scala 380:15:@42389.4]
  assign io_loadHead = head; // @[LoadQueue.scala 379:15:@42388.4]
  assign io_loadEmpty = _T_98323 & _T_98285; // @[LoadQueue.scala 371:16:@42387.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[LoadQueue.scala 382:19:@42406.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[LoadQueue.scala 382:19:@42407.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[LoadQueue.scala 382:19:@42408.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[LoadQueue.scala 382:19:@42409.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[LoadQueue.scala 382:19:@42410.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[LoadQueue.scala 382:19:@42411.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[LoadQueue.scala 382:19:@42412.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[LoadQueue.scala 382:19:@42413.4]
  assign io_loadAddrDone_8 = addrKnown_8; // @[LoadQueue.scala 382:19:@42414.4]
  assign io_loadAddrDone_9 = addrKnown_9; // @[LoadQueue.scala 382:19:@42415.4]
  assign io_loadAddrDone_10 = addrKnown_10; // @[LoadQueue.scala 382:19:@42416.4]
  assign io_loadAddrDone_11 = addrKnown_11; // @[LoadQueue.scala 382:19:@42417.4]
  assign io_loadAddrDone_12 = addrKnown_12; // @[LoadQueue.scala 382:19:@42418.4]
  assign io_loadAddrDone_13 = addrKnown_13; // @[LoadQueue.scala 382:19:@42419.4]
  assign io_loadAddrDone_14 = addrKnown_14; // @[LoadQueue.scala 382:19:@42420.4]
  assign io_loadAddrDone_15 = addrKnown_15; // @[LoadQueue.scala 382:19:@42421.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[LoadQueue.scala 383:19:@42422.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[LoadQueue.scala 383:19:@42423.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[LoadQueue.scala 383:19:@42424.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[LoadQueue.scala 383:19:@42425.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[LoadQueue.scala 383:19:@42426.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[LoadQueue.scala 383:19:@42427.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[LoadQueue.scala 383:19:@42428.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[LoadQueue.scala 383:19:@42429.4]
  assign io_loadDataDone_8 = dataKnown_8; // @[LoadQueue.scala 383:19:@42430.4]
  assign io_loadDataDone_9 = dataKnown_9; // @[LoadQueue.scala 383:19:@42431.4]
  assign io_loadDataDone_10 = dataKnown_10; // @[LoadQueue.scala 383:19:@42432.4]
  assign io_loadDataDone_11 = dataKnown_11; // @[LoadQueue.scala 383:19:@42433.4]
  assign io_loadDataDone_12 = dataKnown_12; // @[LoadQueue.scala 383:19:@42434.4]
  assign io_loadDataDone_13 = dataKnown_13; // @[LoadQueue.scala 383:19:@42435.4]
  assign io_loadDataDone_14 = dataKnown_14; // @[LoadQueue.scala 383:19:@42436.4]
  assign io_loadDataDone_15 = dataKnown_15; // @[LoadQueue.scala 383:19:@42437.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[LoadQueue.scala 381:20:@42390.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[LoadQueue.scala 381:20:@42391.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[LoadQueue.scala 381:20:@42392.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[LoadQueue.scala 381:20:@42393.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[LoadQueue.scala 381:20:@42394.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[LoadQueue.scala 381:20:@42395.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[LoadQueue.scala 381:20:@42396.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[LoadQueue.scala 381:20:@42397.4]
  assign io_loadAddrQueue_8 = addrQ_8; // @[LoadQueue.scala 381:20:@42398.4]
  assign io_loadAddrQueue_9 = addrQ_9; // @[LoadQueue.scala 381:20:@42399.4]
  assign io_loadAddrQueue_10 = addrQ_10; // @[LoadQueue.scala 381:20:@42400.4]
  assign io_loadAddrQueue_11 = addrQ_11; // @[LoadQueue.scala 381:20:@42401.4]
  assign io_loadAddrQueue_12 = addrQ_12; // @[LoadQueue.scala 381:20:@42402.4]
  assign io_loadAddrQueue_13 = addrQ_13; // @[LoadQueue.scala 381:20:@42403.4]
  assign io_loadAddrQueue_14 = addrQ_14; // @[LoadQueue.scala 381:20:@42404.4]
  assign io_loadAddrQueue_15 = addrQ_15; // @[LoadQueue.scala 381:20:@42405.4]
  assign io_loadPorts_0_valid = _T_98182 | _T_98038; // @[LoadQueue.scala 350:38:@42301.6 LoadQueue.scala 353:38:@42305.6]
  assign io_loadPorts_0_bits = _T_98183 ? _GEN_2225 : 32'h0; // @[LoadQueue.scala 349:37:@42300.6 LoadQueue.scala 352:37:@42304.6]
  assign io_loadAddrToMem = _T_93610 ? _GEN_2047 : 32'h0; // @[LoadQueue.scala 248:24:@39139.6 LoadQueue.scala 251:24:@39143.6]
  assign io_loadEnableToMem = _T_93609 | loadRequest_15; // @[LoadQueue.scala 246:22:@39106.4 LoadQueue.scala 249:26:@39140.6 LoadQueue.scala 252:26:@39144.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  loadCompleted_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  loadCompleted_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  loadCompleted_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  loadCompleted_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  loadCompleted_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  loadCompleted_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  loadCompleted_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  loadCompleted_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  bypassInitiated_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  bypassInitiated_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  bypassInitiated_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  bypassInitiated_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  bypassInitiated_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  bypassInitiated_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  bypassInitiated_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  bypassInitiated_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  checkBits_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  checkBits_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  checkBits_2 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  checkBits_3 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  checkBits_4 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  checkBits_5 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  checkBits_6 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  checkBits_7 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  checkBits_8 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  checkBits_9 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  checkBits_10 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  checkBits_11 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  checkBits_12 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  checkBits_13 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  checkBits_14 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  checkBits_15 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  previousStoreHead = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  conflictPReg_0_8 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  conflictPReg_0_9 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  conflictPReg_0_10 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  conflictPReg_0_11 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  conflictPReg_0_12 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  conflictPReg_0_13 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  conflictPReg_0_14 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  conflictPReg_0_15 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  conflictPReg_1_8 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  conflictPReg_1_9 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  conflictPReg_1_10 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  conflictPReg_1_11 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  conflictPReg_1_12 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  conflictPReg_1_13 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  conflictPReg_1_14 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  conflictPReg_1_15 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  conflictPReg_2_8 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  conflictPReg_2_9 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  conflictPReg_2_10 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  conflictPReg_2_11 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  conflictPReg_2_12 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  conflictPReg_2_13 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  conflictPReg_2_14 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  conflictPReg_2_15 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  conflictPReg_3_8 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  conflictPReg_3_9 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  conflictPReg_3_10 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  conflictPReg_3_11 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  conflictPReg_3_12 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  conflictPReg_3_13 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  conflictPReg_3_14 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  conflictPReg_3_15 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  conflictPReg_4_8 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  conflictPReg_4_9 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  conflictPReg_4_10 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  conflictPReg_4_11 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  conflictPReg_4_12 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  conflictPReg_4_13 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  conflictPReg_4_14 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  conflictPReg_4_15 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  conflictPReg_5_8 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  conflictPReg_5_9 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  conflictPReg_5_10 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  conflictPReg_5_11 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  conflictPReg_5_12 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  conflictPReg_5_13 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  conflictPReg_5_14 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  conflictPReg_5_15 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  conflictPReg_6_8 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  conflictPReg_6_9 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  conflictPReg_6_10 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  conflictPReg_6_11 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  conflictPReg_6_12 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  conflictPReg_6_13 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  conflictPReg_6_14 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  conflictPReg_6_15 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  conflictPReg_7_8 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  conflictPReg_7_9 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  conflictPReg_7_10 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  conflictPReg_7_11 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  conflictPReg_7_12 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  conflictPReg_7_13 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  conflictPReg_7_14 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  conflictPReg_7_15 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  conflictPReg_8_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  conflictPReg_8_1 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  conflictPReg_8_2 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  conflictPReg_8_3 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  conflictPReg_8_4 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  conflictPReg_8_5 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  conflictPReg_8_6 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  conflictPReg_8_7 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  conflictPReg_8_8 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  conflictPReg_8_9 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  conflictPReg_8_10 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  conflictPReg_8_11 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  conflictPReg_8_12 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  conflictPReg_8_13 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  conflictPReg_8_14 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  conflictPReg_8_15 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  conflictPReg_9_0 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  conflictPReg_9_1 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  conflictPReg_9_2 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  conflictPReg_9_3 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  conflictPReg_9_4 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  conflictPReg_9_5 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  conflictPReg_9_6 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  conflictPReg_9_7 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  conflictPReg_9_8 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  conflictPReg_9_9 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  conflictPReg_9_10 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  conflictPReg_9_11 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  conflictPReg_9_12 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  conflictPReg_9_13 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  conflictPReg_9_14 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  conflictPReg_9_15 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  conflictPReg_10_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  conflictPReg_10_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  conflictPReg_10_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  conflictPReg_10_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  conflictPReg_10_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  conflictPReg_10_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  conflictPReg_10_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  conflictPReg_10_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  conflictPReg_10_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  conflictPReg_10_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  conflictPReg_10_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  conflictPReg_10_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  conflictPReg_10_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  conflictPReg_10_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  conflictPReg_10_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  conflictPReg_10_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  conflictPReg_11_0 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  conflictPReg_11_1 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  conflictPReg_11_2 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  conflictPReg_11_3 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  conflictPReg_11_4 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  conflictPReg_11_5 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  conflictPReg_11_6 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  conflictPReg_11_7 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  conflictPReg_11_8 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  conflictPReg_11_9 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  conflictPReg_11_10 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  conflictPReg_11_11 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  conflictPReg_11_12 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  conflictPReg_11_13 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  conflictPReg_11_14 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  conflictPReg_11_15 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  conflictPReg_12_0 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  conflictPReg_12_1 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  conflictPReg_12_2 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  conflictPReg_12_3 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  conflictPReg_12_4 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  conflictPReg_12_5 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  conflictPReg_12_6 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  conflictPReg_12_7 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  conflictPReg_12_8 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  conflictPReg_12_9 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  conflictPReg_12_10 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  conflictPReg_12_11 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  conflictPReg_12_12 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  conflictPReg_12_13 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  conflictPReg_12_14 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  conflictPReg_12_15 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  conflictPReg_13_0 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  conflictPReg_13_1 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  conflictPReg_13_2 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  conflictPReg_13_3 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  conflictPReg_13_4 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  conflictPReg_13_5 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  conflictPReg_13_6 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  conflictPReg_13_7 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  conflictPReg_13_8 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  conflictPReg_13_9 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  conflictPReg_13_10 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  conflictPReg_13_11 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  conflictPReg_13_12 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  conflictPReg_13_13 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  conflictPReg_13_14 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  conflictPReg_13_15 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  conflictPReg_14_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  conflictPReg_14_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  conflictPReg_14_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  conflictPReg_14_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  conflictPReg_14_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  conflictPReg_14_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  conflictPReg_14_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  conflictPReg_14_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  conflictPReg_14_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  conflictPReg_14_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  conflictPReg_14_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  conflictPReg_14_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  conflictPReg_14_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  conflictPReg_14_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  conflictPReg_14_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  conflictPReg_14_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  conflictPReg_15_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  conflictPReg_15_1 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  conflictPReg_15_2 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  conflictPReg_15_3 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  conflictPReg_15_4 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  conflictPReg_15_5 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  conflictPReg_15_6 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  conflictPReg_15_7 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  conflictPReg_15_8 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  conflictPReg_15_9 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  conflictPReg_15_10 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  conflictPReg_15_11 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  conflictPReg_15_12 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  conflictPReg_15_13 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  conflictPReg_15_14 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  conflictPReg_15_15 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_8 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_9 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_10 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_11 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_12 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_13 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_14 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_15 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_8 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_9 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_10 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_11 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_12 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_13 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_14 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_15 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_8 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_9 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_10 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_11 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_12 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_13 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_14 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_15 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_8 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_9 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_10 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_11 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_12 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_13 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_14 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_15 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_8 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_9 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_10 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_11 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_12 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_13 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_14 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_15 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_8 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_9 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_10 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_11 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_12 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_13 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_14 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_15 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_8 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_9 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_10 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_11 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_12 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_13 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_14 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_15 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_8 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_9 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_10 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_11 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_12 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_13 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_14 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_15 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_0 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_1 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_2 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_3 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_4 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_5 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_6 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_7 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_8 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_9 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_10 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_11 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_12 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_13 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_14 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_15 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_0 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_1 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_2 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_3 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_4 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_5 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_6 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_7 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_8 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_9 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_10 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_11 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_12 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_13 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_14 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_15 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_0 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_1 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_2 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_3 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_4 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_5 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_6 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_7 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_8 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_9 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_10 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_11 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_12 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_13 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_14 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_15 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_0 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_1 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_2 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_3 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_4 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_5 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_6 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_7 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_8 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_9 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_10 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_11 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_12 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_13 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_14 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_15 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_0 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_1 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_2 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_3 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_4 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_5 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_6 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_7 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_8 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_9 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_10 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_11 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_12 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_13 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_14 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_15 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_0 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_1 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_2 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_3 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_4 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_5 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_6 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_7 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_8 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_9 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_10 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_11 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_12 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_13 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_14 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_15 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_0 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_1 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_2 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_3 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_4 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_5 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_6 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_7 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_8 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_9 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_10 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_11 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_12 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_13 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_14 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_15 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_0 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_1 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_2 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_3 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_4 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_5 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_6 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_7 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_8 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_9 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_10 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_11 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_12 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_13 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_14 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_15 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_8 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_9 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_10 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_11 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_12 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_13 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_14 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_15 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  shiftedStoreDataQPreg_8 = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  shiftedStoreDataQPreg_9 = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  shiftedStoreDataQPreg_10 = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  shiftedStoreDataQPreg_11 = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  shiftedStoreDataQPreg_12 = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  shiftedStoreDataQPreg_13 = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  shiftedStoreDataQPreg_14 = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  shiftedStoreDataQPreg_15 = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  addrKnownPReg_8 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  addrKnownPReg_9 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  addrKnownPReg_10 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  addrKnownPReg_11 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  addrKnownPReg_12 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  addrKnownPReg_13 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  addrKnownPReg_14 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  addrKnownPReg_15 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  dataKnownPReg_8 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  dataKnownPReg_9 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  dataKnownPReg_10 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  dataKnownPReg_11 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  dataKnownPReg_12 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  dataKnownPReg_13 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  dataKnownPReg_14 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  dataKnownPReg_15 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  prevPriorityRequest_15 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  prevPriorityRequest_14 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  prevPriorityRequest_13 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  prevPriorityRequest_12 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  prevPriorityRequest_11 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  prevPriorityRequest_10 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  prevPriorityRequest_9 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  prevPriorityRequest_8 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  prevPriorityRequest_7 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  prevPriorityRequest_6 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  prevPriorityRequest_5 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  prevPriorityRequest_4 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  prevPriorityRequest_3 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  prevPriorityRequest_2 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  prevPriorityRequest_1 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  prevPriorityRequest_0 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_2260[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_2261[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1924) begin
          offsetQ_0 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1924) begin
            offsetQ_0 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1924) begin
              offsetQ_0 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1924) begin
                offsetQ_0 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1924) begin
                  offsetQ_0 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1924) begin
                    offsetQ_0 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1924) begin
                      offsetQ_0 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1924) begin
                        offsetQ_0 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1924) begin
                          offsetQ_0 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1924) begin
                            offsetQ_0 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1924) begin
                              offsetQ_0 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1924) begin
                                offsetQ_0 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1924) begin
                                  offsetQ_0 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1924) begin
                                    offsetQ_0 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1924) begin
                                      offsetQ_0 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1942) begin
          offsetQ_1 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1942) begin
            offsetQ_1 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1942) begin
              offsetQ_1 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1942) begin
                offsetQ_1 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1942) begin
                  offsetQ_1 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1942) begin
                    offsetQ_1 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1942) begin
                      offsetQ_1 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1942) begin
                        offsetQ_1 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1942) begin
                          offsetQ_1 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1942) begin
                            offsetQ_1 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1942) begin
                              offsetQ_1 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1942) begin
                                offsetQ_1 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1942) begin
                                  offsetQ_1 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1942) begin
                                    offsetQ_1 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1942) begin
                                      offsetQ_1 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1960) begin
          offsetQ_2 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1960) begin
            offsetQ_2 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1960) begin
              offsetQ_2 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1960) begin
                offsetQ_2 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1960) begin
                  offsetQ_2 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1960) begin
                    offsetQ_2 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1960) begin
                      offsetQ_2 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1960) begin
                        offsetQ_2 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1960) begin
                          offsetQ_2 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1960) begin
                            offsetQ_2 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1960) begin
                              offsetQ_2 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1960) begin
                                offsetQ_2 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1960) begin
                                  offsetQ_2 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1960) begin
                                    offsetQ_2 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1960) begin
                                      offsetQ_2 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1978) begin
          offsetQ_3 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1978) begin
            offsetQ_3 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1978) begin
              offsetQ_3 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1978) begin
                offsetQ_3 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1978) begin
                  offsetQ_3 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1978) begin
                    offsetQ_3 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1978) begin
                      offsetQ_3 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1978) begin
                        offsetQ_3 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1978) begin
                          offsetQ_3 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1978) begin
                            offsetQ_3 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1978) begin
                              offsetQ_3 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1978) begin
                                offsetQ_3 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1978) begin
                                  offsetQ_3 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1978) begin
                                    offsetQ_3 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1978) begin
                                      offsetQ_3 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1996) begin
          offsetQ_4 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1996) begin
            offsetQ_4 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1996) begin
              offsetQ_4 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1996) begin
                offsetQ_4 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1996) begin
                  offsetQ_4 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1996) begin
                    offsetQ_4 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1996) begin
                      offsetQ_4 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1996) begin
                        offsetQ_4 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1996) begin
                          offsetQ_4 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1996) begin
                            offsetQ_4 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1996) begin
                              offsetQ_4 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1996) begin
                                offsetQ_4 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1996) begin
                                  offsetQ_4 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1996) begin
                                    offsetQ_4 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1996) begin
                                      offsetQ_4 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_2014) begin
          offsetQ_5 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2014) begin
            offsetQ_5 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2014) begin
              offsetQ_5 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2014) begin
                offsetQ_5 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2014) begin
                  offsetQ_5 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2014) begin
                    offsetQ_5 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2014) begin
                      offsetQ_5 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2014) begin
                        offsetQ_5 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2014) begin
                          offsetQ_5 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2014) begin
                            offsetQ_5 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2014) begin
                              offsetQ_5 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2014) begin
                                offsetQ_5 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2014) begin
                                  offsetQ_5 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2014) begin
                                    offsetQ_5 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2014) begin
                                      offsetQ_5 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_2032) begin
          offsetQ_6 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2032) begin
            offsetQ_6 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2032) begin
              offsetQ_6 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2032) begin
                offsetQ_6 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2032) begin
                  offsetQ_6 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2032) begin
                    offsetQ_6 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2032) begin
                      offsetQ_6 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2032) begin
                        offsetQ_6 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2032) begin
                          offsetQ_6 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2032) begin
                            offsetQ_6 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2032) begin
                              offsetQ_6 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2032) begin
                                offsetQ_6 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2032) begin
                                  offsetQ_6 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2032) begin
                                    offsetQ_6 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2032) begin
                                      offsetQ_6 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_2050) begin
          offsetQ_7 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2050) begin
            offsetQ_7 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2050) begin
              offsetQ_7 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2050) begin
                offsetQ_7 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2050) begin
                  offsetQ_7 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2050) begin
                    offsetQ_7 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2050) begin
                      offsetQ_7 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2050) begin
                        offsetQ_7 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2050) begin
                          offsetQ_7 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2050) begin
                            offsetQ_7 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2050) begin
                              offsetQ_7 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2050) begin
                                offsetQ_7 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2050) begin
                                  offsetQ_7 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2050) begin
                                    offsetQ_7 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2050) begin
                                      offsetQ_7 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_2068) begin
          offsetQ_8 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2068) begin
            offsetQ_8 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2068) begin
              offsetQ_8 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2068) begin
                offsetQ_8 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2068) begin
                  offsetQ_8 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2068) begin
                    offsetQ_8 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2068) begin
                      offsetQ_8 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2068) begin
                        offsetQ_8 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2068) begin
                          offsetQ_8 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2068) begin
                            offsetQ_8 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2068) begin
                              offsetQ_8 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2068) begin
                                offsetQ_8 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2068) begin
                                  offsetQ_8 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2068) begin
                                    offsetQ_8 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2068) begin
                                      offsetQ_8 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_2086) begin
          offsetQ_9 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2086) begin
            offsetQ_9 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2086) begin
              offsetQ_9 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2086) begin
                offsetQ_9 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2086) begin
                  offsetQ_9 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2086) begin
                    offsetQ_9 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2086) begin
                      offsetQ_9 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2086) begin
                        offsetQ_9 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2086) begin
                          offsetQ_9 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2086) begin
                            offsetQ_9 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2086) begin
                              offsetQ_9 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2086) begin
                                offsetQ_9 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2086) begin
                                  offsetQ_9 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2086) begin
                                    offsetQ_9 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2086) begin
                                      offsetQ_9 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_2104) begin
          offsetQ_10 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2104) begin
            offsetQ_10 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2104) begin
              offsetQ_10 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2104) begin
                offsetQ_10 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2104) begin
                  offsetQ_10 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2104) begin
                    offsetQ_10 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2104) begin
                      offsetQ_10 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2104) begin
                        offsetQ_10 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2104) begin
                          offsetQ_10 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2104) begin
                            offsetQ_10 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2104) begin
                              offsetQ_10 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2104) begin
                                offsetQ_10 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2104) begin
                                  offsetQ_10 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2104) begin
                                    offsetQ_10 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2104) begin
                                      offsetQ_10 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2122) begin
          offsetQ_11 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2122) begin
            offsetQ_11 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2122) begin
              offsetQ_11 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2122) begin
                offsetQ_11 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2122) begin
                  offsetQ_11 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2122) begin
                    offsetQ_11 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2122) begin
                      offsetQ_11 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2122) begin
                        offsetQ_11 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2122) begin
                          offsetQ_11 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2122) begin
                            offsetQ_11 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2122) begin
                              offsetQ_11 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2122) begin
                                offsetQ_11 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2122) begin
                                  offsetQ_11 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2122) begin
                                    offsetQ_11 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2122) begin
                                      offsetQ_11 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2140) begin
          offsetQ_12 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2140) begin
            offsetQ_12 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2140) begin
              offsetQ_12 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2140) begin
                offsetQ_12 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2140) begin
                  offsetQ_12 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2140) begin
                    offsetQ_12 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2140) begin
                      offsetQ_12 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2140) begin
                        offsetQ_12 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2140) begin
                          offsetQ_12 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2140) begin
                            offsetQ_12 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2140) begin
                              offsetQ_12 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2140) begin
                                offsetQ_12 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2140) begin
                                  offsetQ_12 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2140) begin
                                    offsetQ_12 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2140) begin
                                      offsetQ_12 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2158) begin
          offsetQ_13 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2158) begin
            offsetQ_13 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2158) begin
              offsetQ_13 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2158) begin
                offsetQ_13 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2158) begin
                  offsetQ_13 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2158) begin
                    offsetQ_13 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2158) begin
                      offsetQ_13 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2158) begin
                        offsetQ_13 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2158) begin
                          offsetQ_13 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2158) begin
                            offsetQ_13 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2158) begin
                              offsetQ_13 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2158) begin
                                offsetQ_13 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2158) begin
                                  offsetQ_13 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2158) begin
                                    offsetQ_13 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2158) begin
                                      offsetQ_13 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2176) begin
          offsetQ_14 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2176) begin
            offsetQ_14 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2176) begin
              offsetQ_14 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2176) begin
                offsetQ_14 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2176) begin
                  offsetQ_14 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2176) begin
                    offsetQ_14 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2176) begin
                      offsetQ_14 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2176) begin
                        offsetQ_14 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2176) begin
                          offsetQ_14 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2176) begin
                            offsetQ_14 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2176) begin
                              offsetQ_14 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2176) begin
                                offsetQ_14 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2176) begin
                                  offsetQ_14 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2176) begin
                                    offsetQ_14 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2176) begin
                                      offsetQ_14 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2194) begin
          offsetQ_15 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2194) begin
            offsetQ_15 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2194) begin
              offsetQ_15 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2194) begin
                offsetQ_15 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2194) begin
                  offsetQ_15 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2194) begin
                    offsetQ_15 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2194) begin
                      offsetQ_15 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2194) begin
                        offsetQ_15 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2194) begin
                          offsetQ_15 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2194) begin
                            offsetQ_15 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2194) begin
                              offsetQ_15 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2194) begin
                                offsetQ_15 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2194) begin
                                  offsetQ_15 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2194) begin
                                    offsetQ_15 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2194) begin
                                      offsetQ_15 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_97565) begin
          addrQ_0 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_97580) begin
          addrQ_1 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_97595) begin
          addrQ_2 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_97610) begin
          addrQ_3 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_97625) begin
          addrQ_4 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_97640) begin
          addrQ_5 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_97655) begin
          addrQ_6 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_97670) begin
          addrQ_7 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_97685) begin
          addrQ_8 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_97700) begin
          addrQ_9 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_97715) begin
          addrQ_10 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_97730) begin
          addrQ_11 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_97745) begin
          addrQ_12 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_97760) begin
          addrQ_13 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_97775) begin
          addrQ_14 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_97790) begin
          addrQ_15 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_88298) begin
          if (4'hf == _T_88281) begin
            dataQ_0 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88281) begin
              dataQ_0 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88281) begin
                dataQ_0 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88281) begin
                  dataQ_0 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88281) begin
                    dataQ_0 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88281) begin
                      dataQ_0 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88281) begin
                        dataQ_0 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88281) begin
                          dataQ_0 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88281) begin
                            dataQ_0 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88281) begin
                              dataQ_0 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88281) begin
                                dataQ_0 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88281) begin
                                  dataQ_0 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88281) begin
                                    dataQ_0 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88281) begin
                                      dataQ_0 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88281) begin
                                        dataQ_0 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_0 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_0) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_88434) begin
          if (4'hf == _T_88417) begin
            dataQ_1 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88417) begin
              dataQ_1 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88417) begin
                dataQ_1 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88417) begin
                  dataQ_1 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88417) begin
                    dataQ_1 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88417) begin
                      dataQ_1 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88417) begin
                        dataQ_1 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88417) begin
                          dataQ_1 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88417) begin
                            dataQ_1 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88417) begin
                              dataQ_1 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88417) begin
                                dataQ_1 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88417) begin
                                  dataQ_1 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88417) begin
                                    dataQ_1 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88417) begin
                                      dataQ_1 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88417) begin
                                        dataQ_1 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_1 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_1) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_88570) begin
          if (4'hf == _T_88553) begin
            dataQ_2 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88553) begin
              dataQ_2 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88553) begin
                dataQ_2 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88553) begin
                  dataQ_2 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88553) begin
                    dataQ_2 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88553) begin
                      dataQ_2 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88553) begin
                        dataQ_2 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88553) begin
                          dataQ_2 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88553) begin
                            dataQ_2 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88553) begin
                              dataQ_2 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88553) begin
                                dataQ_2 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88553) begin
                                  dataQ_2 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88553) begin
                                    dataQ_2 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88553) begin
                                      dataQ_2 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88553) begin
                                        dataQ_2 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_2 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_2) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_88706) begin
          if (4'hf == _T_88689) begin
            dataQ_3 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88689) begin
              dataQ_3 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88689) begin
                dataQ_3 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88689) begin
                  dataQ_3 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88689) begin
                    dataQ_3 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88689) begin
                      dataQ_3 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88689) begin
                        dataQ_3 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88689) begin
                          dataQ_3 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88689) begin
                            dataQ_3 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88689) begin
                              dataQ_3 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88689) begin
                                dataQ_3 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88689) begin
                                  dataQ_3 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88689) begin
                                    dataQ_3 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88689) begin
                                      dataQ_3 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88689) begin
                                        dataQ_3 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_3 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_3) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_88842) begin
          if (4'hf == _T_88825) begin
            dataQ_4 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88825) begin
              dataQ_4 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88825) begin
                dataQ_4 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88825) begin
                  dataQ_4 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88825) begin
                    dataQ_4 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88825) begin
                      dataQ_4 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88825) begin
                        dataQ_4 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88825) begin
                          dataQ_4 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88825) begin
                            dataQ_4 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88825) begin
                              dataQ_4 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88825) begin
                                dataQ_4 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88825) begin
                                  dataQ_4 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88825) begin
                                    dataQ_4 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88825) begin
                                      dataQ_4 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88825) begin
                                        dataQ_4 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_4 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_4) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_88978) begin
          if (4'hf == _T_88961) begin
            dataQ_5 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88961) begin
              dataQ_5 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88961) begin
                dataQ_5 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88961) begin
                  dataQ_5 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88961) begin
                    dataQ_5 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88961) begin
                      dataQ_5 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88961) begin
                        dataQ_5 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88961) begin
                          dataQ_5 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88961) begin
                            dataQ_5 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88961) begin
                              dataQ_5 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88961) begin
                                dataQ_5 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88961) begin
                                  dataQ_5 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88961) begin
                                    dataQ_5 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88961) begin
                                      dataQ_5 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88961) begin
                                        dataQ_5 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_5 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_5) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_89114) begin
          if (4'hf == _T_89097) begin
            dataQ_6 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89097) begin
              dataQ_6 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89097) begin
                dataQ_6 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89097) begin
                  dataQ_6 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89097) begin
                    dataQ_6 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89097) begin
                      dataQ_6 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89097) begin
                        dataQ_6 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89097) begin
                          dataQ_6 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89097) begin
                            dataQ_6 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89097) begin
                              dataQ_6 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89097) begin
                                dataQ_6 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89097) begin
                                  dataQ_6 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89097) begin
                                    dataQ_6 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89097) begin
                                      dataQ_6 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89097) begin
                                        dataQ_6 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_6 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_6) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_89250) begin
          if (4'hf == _T_89233) begin
            dataQ_7 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89233) begin
              dataQ_7 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89233) begin
                dataQ_7 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89233) begin
                  dataQ_7 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89233) begin
                    dataQ_7 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89233) begin
                      dataQ_7 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89233) begin
                        dataQ_7 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89233) begin
                          dataQ_7 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89233) begin
                            dataQ_7 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89233) begin
                              dataQ_7 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89233) begin
                                dataQ_7 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89233) begin
                                  dataQ_7 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89233) begin
                                    dataQ_7 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89233) begin
                                      dataQ_7 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89233) begin
                                        dataQ_7 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_7 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_7) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (bypassRequest_8) begin
        if (_T_89386) begin
          if (4'hf == _T_89369) begin
            dataQ_8 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89369) begin
              dataQ_8 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89369) begin
                dataQ_8 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89369) begin
                  dataQ_8 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89369) begin
                    dataQ_8 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89369) begin
                      dataQ_8 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89369) begin
                        dataQ_8 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89369) begin
                          dataQ_8 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89369) begin
                            dataQ_8 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89369) begin
                              dataQ_8 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89369) begin
                                dataQ_8 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89369) begin
                                  dataQ_8 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89369) begin
                                    dataQ_8 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89369) begin
                                      dataQ_8 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89369) begin
                                        dataQ_8 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_8 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_8 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_8) begin
          dataQ_8 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (bypassRequest_9) begin
        if (_T_89522) begin
          if (4'hf == _T_89505) begin
            dataQ_9 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89505) begin
              dataQ_9 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89505) begin
                dataQ_9 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89505) begin
                  dataQ_9 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89505) begin
                    dataQ_9 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89505) begin
                      dataQ_9 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89505) begin
                        dataQ_9 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89505) begin
                          dataQ_9 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89505) begin
                            dataQ_9 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89505) begin
                              dataQ_9 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89505) begin
                                dataQ_9 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89505) begin
                                  dataQ_9 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89505) begin
                                    dataQ_9 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89505) begin
                                      dataQ_9 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89505) begin
                                        dataQ_9 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_9 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_9 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_9) begin
          dataQ_9 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (bypassRequest_10) begin
        if (_T_89658) begin
          if (4'hf == _T_89641) begin
            dataQ_10 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89641) begin
              dataQ_10 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89641) begin
                dataQ_10 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89641) begin
                  dataQ_10 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89641) begin
                    dataQ_10 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89641) begin
                      dataQ_10 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89641) begin
                        dataQ_10 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89641) begin
                          dataQ_10 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89641) begin
                            dataQ_10 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89641) begin
                              dataQ_10 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89641) begin
                                dataQ_10 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89641) begin
                                  dataQ_10 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89641) begin
                                    dataQ_10 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89641) begin
                                      dataQ_10 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89641) begin
                                        dataQ_10 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_10 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_10 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_10) begin
          dataQ_10 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (bypassRequest_11) begin
        if (_T_89794) begin
          if (4'hf == _T_89777) begin
            dataQ_11 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89777) begin
              dataQ_11 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89777) begin
                dataQ_11 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89777) begin
                  dataQ_11 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89777) begin
                    dataQ_11 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89777) begin
                      dataQ_11 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89777) begin
                        dataQ_11 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89777) begin
                          dataQ_11 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89777) begin
                            dataQ_11 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89777) begin
                              dataQ_11 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89777) begin
                                dataQ_11 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89777) begin
                                  dataQ_11 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89777) begin
                                    dataQ_11 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89777) begin
                                      dataQ_11 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89777) begin
                                        dataQ_11 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_11 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_11 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_11) begin
          dataQ_11 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (bypassRequest_12) begin
        if (_T_89930) begin
          if (4'hf == _T_89913) begin
            dataQ_12 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89913) begin
              dataQ_12 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89913) begin
                dataQ_12 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89913) begin
                  dataQ_12 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89913) begin
                    dataQ_12 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89913) begin
                      dataQ_12 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89913) begin
                        dataQ_12 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89913) begin
                          dataQ_12 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89913) begin
                            dataQ_12 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89913) begin
                              dataQ_12 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89913) begin
                                dataQ_12 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89913) begin
                                  dataQ_12 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89913) begin
                                    dataQ_12 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89913) begin
                                      dataQ_12 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89913) begin
                                        dataQ_12 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_12 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_12 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_12) begin
          dataQ_12 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (bypassRequest_13) begin
        if (_T_90066) begin
          if (4'hf == _T_90049) begin
            dataQ_13 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90049) begin
              dataQ_13 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90049) begin
                dataQ_13 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90049) begin
                  dataQ_13 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90049) begin
                    dataQ_13 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90049) begin
                      dataQ_13 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90049) begin
                        dataQ_13 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90049) begin
                          dataQ_13 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90049) begin
                            dataQ_13 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90049) begin
                              dataQ_13 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90049) begin
                                dataQ_13 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90049) begin
                                  dataQ_13 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90049) begin
                                    dataQ_13 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90049) begin
                                      dataQ_13 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90049) begin
                                        dataQ_13 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_13 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_13 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_13) begin
          dataQ_13 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (bypassRequest_14) begin
        if (_T_90202) begin
          if (4'hf == _T_90185) begin
            dataQ_14 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90185) begin
              dataQ_14 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90185) begin
                dataQ_14 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90185) begin
                  dataQ_14 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90185) begin
                    dataQ_14 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90185) begin
                      dataQ_14 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90185) begin
                        dataQ_14 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90185) begin
                          dataQ_14 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90185) begin
                            dataQ_14 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90185) begin
                              dataQ_14 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90185) begin
                                dataQ_14 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90185) begin
                                  dataQ_14 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90185) begin
                                    dataQ_14 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90185) begin
                                      dataQ_14 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90185) begin
                                        dataQ_14 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_14 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_14 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_14) begin
          dataQ_14 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (bypassRequest_15) begin
        if (_T_90338) begin
          if (4'hf == _T_90321) begin
            dataQ_15 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90321) begin
              dataQ_15 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90321) begin
                dataQ_15 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90321) begin
                  dataQ_15 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90321) begin
                    dataQ_15 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90321) begin
                      dataQ_15 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90321) begin
                        dataQ_15 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90321) begin
                          dataQ_15 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90321) begin
                            dataQ_15 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90321) begin
                              dataQ_15 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90321) begin
                                dataQ_15 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90321) begin
                                  dataQ_15 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90321) begin
                                    dataQ_15 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90321) begin
                                      dataQ_15 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90321) begin
                                        dataQ_15 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_15 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_15 <= 32'h0;
        end
      end else begin
        if (prevPriorityRequest_15) begin
          dataQ_15 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_97565) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_97580) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_97595) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_97610) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_97625) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_97640) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_97655) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_97670) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_97685) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_97700) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_97715) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_97730) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_97745) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_97760) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_97775) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_97790) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_93649) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_93652) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_93655) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_93658) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_93661) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_93664) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_93667) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_93670) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_93673) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_93676) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_93679) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_93682) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_93685) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_93688) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_93691) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_93694) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        loadCompleted_8 <= 1'h0;
      end else begin
        if (loadCompleting_8) begin
          loadCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        loadCompleted_9 <= 1'h0;
      end else begin
        if (loadCompleting_9) begin
          loadCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        loadCompleted_10 <= 1'h0;
      end else begin
        if (loadCompleting_10) begin
          loadCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        loadCompleted_11 <= 1'h0;
      end else begin
        if (loadCompleting_11) begin
          loadCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        loadCompleted_12 <= 1'h0;
      end else begin
        if (loadCompleting_12) begin
          loadCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        loadCompleted_13 <= 1'h0;
      end else begin
        if (loadCompleting_13) begin
          loadCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        loadCompleted_14 <= 1'h0;
      end else begin
        if (loadCompleting_14) begin
          loadCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        loadCompleted_15 <= 1'h0;
      end else begin
        if (loadCompleting_15) begin
          loadCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1878;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1879;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1880;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1881;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1882;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1883;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1884;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1885;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1886;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1887;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1888;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1889;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1890;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1891;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1892;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1893;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        bypassInitiated_8 <= 1'h0;
      end else begin
        if (bypassRequest_8) begin
          bypassInitiated_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        bypassInitiated_9 <= 1'h0;
      end else begin
        if (bypassRequest_9) begin
          bypassInitiated_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        bypassInitiated_10 <= 1'h0;
      end else begin
        if (bypassRequest_10) begin
          bypassInitiated_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        bypassInitiated_11 <= 1'h0;
      end else begin
        if (bypassRequest_11) begin
          bypassInitiated_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        bypassInitiated_12 <= 1'h0;
      end else begin
        if (bypassRequest_12) begin
          bypassInitiated_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        bypassInitiated_13 <= 1'h0;
      end else begin
        if (bypassRequest_13) begin
          bypassInitiated_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        bypassInitiated_14 <= 1'h0;
      end else begin
        if (bypassRequest_14) begin
          bypassInitiated_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        bypassInitiated_15 <= 1'h0;
      end else begin
        if (bypassRequest_15) begin
          bypassInitiated_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2221;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2225) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2233) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2251;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2255) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2263) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2281;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2285) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2293) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2311;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2315) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2323) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2341;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2345) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2353) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2371;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2375) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2383) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2401;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2405) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2413) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2431;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2435) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2443) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2461;
      end else begin
        if (io_storeEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2465) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2473) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2491;
      end else begin
        if (io_storeEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2495) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2503) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2521;
      end else begin
        if (io_storeEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2525) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2533) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2551;
      end else begin
        if (io_storeEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2555) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2563) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2581;
      end else begin
        if (io_storeEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2585) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2593) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2611;
      end else begin
        if (io_storeEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2615) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2623) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2641;
      end else begin
        if (io_storeEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2645) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2653) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2671;
      end else begin
        if (io_storeEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2675) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2683) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_18282[0];
    conflictPReg_0_1 <= _T_18282[1];
    conflictPReg_0_2 <= _T_18282[2];
    conflictPReg_0_3 <= _T_18282[3];
    conflictPReg_0_4 <= _T_18282[4];
    conflictPReg_0_5 <= _T_18282[5];
    conflictPReg_0_6 <= _T_18282[6];
    conflictPReg_0_7 <= _T_18282[7];
    conflictPReg_0_8 <= _T_18282[8];
    conflictPReg_0_9 <= _T_18282[9];
    conflictPReg_0_10 <= _T_18282[10];
    conflictPReg_0_11 <= _T_18282[11];
    conflictPReg_0_12 <= _T_18282[12];
    conflictPReg_0_13 <= _T_18282[13];
    conflictPReg_0_14 <= _T_18282[14];
    conflictPReg_0_15 <= _T_18282[15];
    conflictPReg_1_0 <= _T_19140[0];
    conflictPReg_1_1 <= _T_19140[1];
    conflictPReg_1_2 <= _T_19140[2];
    conflictPReg_1_3 <= _T_19140[3];
    conflictPReg_1_4 <= _T_19140[4];
    conflictPReg_1_5 <= _T_19140[5];
    conflictPReg_1_6 <= _T_19140[6];
    conflictPReg_1_7 <= _T_19140[7];
    conflictPReg_1_8 <= _T_19140[8];
    conflictPReg_1_9 <= _T_19140[9];
    conflictPReg_1_10 <= _T_19140[10];
    conflictPReg_1_11 <= _T_19140[11];
    conflictPReg_1_12 <= _T_19140[12];
    conflictPReg_1_13 <= _T_19140[13];
    conflictPReg_1_14 <= _T_19140[14];
    conflictPReg_1_15 <= _T_19140[15];
    conflictPReg_2_0 <= _T_19998[0];
    conflictPReg_2_1 <= _T_19998[1];
    conflictPReg_2_2 <= _T_19998[2];
    conflictPReg_2_3 <= _T_19998[3];
    conflictPReg_2_4 <= _T_19998[4];
    conflictPReg_2_5 <= _T_19998[5];
    conflictPReg_2_6 <= _T_19998[6];
    conflictPReg_2_7 <= _T_19998[7];
    conflictPReg_2_8 <= _T_19998[8];
    conflictPReg_2_9 <= _T_19998[9];
    conflictPReg_2_10 <= _T_19998[10];
    conflictPReg_2_11 <= _T_19998[11];
    conflictPReg_2_12 <= _T_19998[12];
    conflictPReg_2_13 <= _T_19998[13];
    conflictPReg_2_14 <= _T_19998[14];
    conflictPReg_2_15 <= _T_19998[15];
    conflictPReg_3_0 <= _T_20856[0];
    conflictPReg_3_1 <= _T_20856[1];
    conflictPReg_3_2 <= _T_20856[2];
    conflictPReg_3_3 <= _T_20856[3];
    conflictPReg_3_4 <= _T_20856[4];
    conflictPReg_3_5 <= _T_20856[5];
    conflictPReg_3_6 <= _T_20856[6];
    conflictPReg_3_7 <= _T_20856[7];
    conflictPReg_3_8 <= _T_20856[8];
    conflictPReg_3_9 <= _T_20856[9];
    conflictPReg_3_10 <= _T_20856[10];
    conflictPReg_3_11 <= _T_20856[11];
    conflictPReg_3_12 <= _T_20856[12];
    conflictPReg_3_13 <= _T_20856[13];
    conflictPReg_3_14 <= _T_20856[14];
    conflictPReg_3_15 <= _T_20856[15];
    conflictPReg_4_0 <= _T_21714[0];
    conflictPReg_4_1 <= _T_21714[1];
    conflictPReg_4_2 <= _T_21714[2];
    conflictPReg_4_3 <= _T_21714[3];
    conflictPReg_4_4 <= _T_21714[4];
    conflictPReg_4_5 <= _T_21714[5];
    conflictPReg_4_6 <= _T_21714[6];
    conflictPReg_4_7 <= _T_21714[7];
    conflictPReg_4_8 <= _T_21714[8];
    conflictPReg_4_9 <= _T_21714[9];
    conflictPReg_4_10 <= _T_21714[10];
    conflictPReg_4_11 <= _T_21714[11];
    conflictPReg_4_12 <= _T_21714[12];
    conflictPReg_4_13 <= _T_21714[13];
    conflictPReg_4_14 <= _T_21714[14];
    conflictPReg_4_15 <= _T_21714[15];
    conflictPReg_5_0 <= _T_22572[0];
    conflictPReg_5_1 <= _T_22572[1];
    conflictPReg_5_2 <= _T_22572[2];
    conflictPReg_5_3 <= _T_22572[3];
    conflictPReg_5_4 <= _T_22572[4];
    conflictPReg_5_5 <= _T_22572[5];
    conflictPReg_5_6 <= _T_22572[6];
    conflictPReg_5_7 <= _T_22572[7];
    conflictPReg_5_8 <= _T_22572[8];
    conflictPReg_5_9 <= _T_22572[9];
    conflictPReg_5_10 <= _T_22572[10];
    conflictPReg_5_11 <= _T_22572[11];
    conflictPReg_5_12 <= _T_22572[12];
    conflictPReg_5_13 <= _T_22572[13];
    conflictPReg_5_14 <= _T_22572[14];
    conflictPReg_5_15 <= _T_22572[15];
    conflictPReg_6_0 <= _T_23430[0];
    conflictPReg_6_1 <= _T_23430[1];
    conflictPReg_6_2 <= _T_23430[2];
    conflictPReg_6_3 <= _T_23430[3];
    conflictPReg_6_4 <= _T_23430[4];
    conflictPReg_6_5 <= _T_23430[5];
    conflictPReg_6_6 <= _T_23430[6];
    conflictPReg_6_7 <= _T_23430[7];
    conflictPReg_6_8 <= _T_23430[8];
    conflictPReg_6_9 <= _T_23430[9];
    conflictPReg_6_10 <= _T_23430[10];
    conflictPReg_6_11 <= _T_23430[11];
    conflictPReg_6_12 <= _T_23430[12];
    conflictPReg_6_13 <= _T_23430[13];
    conflictPReg_6_14 <= _T_23430[14];
    conflictPReg_6_15 <= _T_23430[15];
    conflictPReg_7_0 <= _T_24288[0];
    conflictPReg_7_1 <= _T_24288[1];
    conflictPReg_7_2 <= _T_24288[2];
    conflictPReg_7_3 <= _T_24288[3];
    conflictPReg_7_4 <= _T_24288[4];
    conflictPReg_7_5 <= _T_24288[5];
    conflictPReg_7_6 <= _T_24288[6];
    conflictPReg_7_7 <= _T_24288[7];
    conflictPReg_7_8 <= _T_24288[8];
    conflictPReg_7_9 <= _T_24288[9];
    conflictPReg_7_10 <= _T_24288[10];
    conflictPReg_7_11 <= _T_24288[11];
    conflictPReg_7_12 <= _T_24288[12];
    conflictPReg_7_13 <= _T_24288[13];
    conflictPReg_7_14 <= _T_24288[14];
    conflictPReg_7_15 <= _T_24288[15];
    conflictPReg_8_0 <= _T_25146[0];
    conflictPReg_8_1 <= _T_25146[1];
    conflictPReg_8_2 <= _T_25146[2];
    conflictPReg_8_3 <= _T_25146[3];
    conflictPReg_8_4 <= _T_25146[4];
    conflictPReg_8_5 <= _T_25146[5];
    conflictPReg_8_6 <= _T_25146[6];
    conflictPReg_8_7 <= _T_25146[7];
    conflictPReg_8_8 <= _T_25146[8];
    conflictPReg_8_9 <= _T_25146[9];
    conflictPReg_8_10 <= _T_25146[10];
    conflictPReg_8_11 <= _T_25146[11];
    conflictPReg_8_12 <= _T_25146[12];
    conflictPReg_8_13 <= _T_25146[13];
    conflictPReg_8_14 <= _T_25146[14];
    conflictPReg_8_15 <= _T_25146[15];
    conflictPReg_9_0 <= _T_26004[0];
    conflictPReg_9_1 <= _T_26004[1];
    conflictPReg_9_2 <= _T_26004[2];
    conflictPReg_9_3 <= _T_26004[3];
    conflictPReg_9_4 <= _T_26004[4];
    conflictPReg_9_5 <= _T_26004[5];
    conflictPReg_9_6 <= _T_26004[6];
    conflictPReg_9_7 <= _T_26004[7];
    conflictPReg_9_8 <= _T_26004[8];
    conflictPReg_9_9 <= _T_26004[9];
    conflictPReg_9_10 <= _T_26004[10];
    conflictPReg_9_11 <= _T_26004[11];
    conflictPReg_9_12 <= _T_26004[12];
    conflictPReg_9_13 <= _T_26004[13];
    conflictPReg_9_14 <= _T_26004[14];
    conflictPReg_9_15 <= _T_26004[15];
    conflictPReg_10_0 <= _T_26862[0];
    conflictPReg_10_1 <= _T_26862[1];
    conflictPReg_10_2 <= _T_26862[2];
    conflictPReg_10_3 <= _T_26862[3];
    conflictPReg_10_4 <= _T_26862[4];
    conflictPReg_10_5 <= _T_26862[5];
    conflictPReg_10_6 <= _T_26862[6];
    conflictPReg_10_7 <= _T_26862[7];
    conflictPReg_10_8 <= _T_26862[8];
    conflictPReg_10_9 <= _T_26862[9];
    conflictPReg_10_10 <= _T_26862[10];
    conflictPReg_10_11 <= _T_26862[11];
    conflictPReg_10_12 <= _T_26862[12];
    conflictPReg_10_13 <= _T_26862[13];
    conflictPReg_10_14 <= _T_26862[14];
    conflictPReg_10_15 <= _T_26862[15];
    conflictPReg_11_0 <= _T_27720[0];
    conflictPReg_11_1 <= _T_27720[1];
    conflictPReg_11_2 <= _T_27720[2];
    conflictPReg_11_3 <= _T_27720[3];
    conflictPReg_11_4 <= _T_27720[4];
    conflictPReg_11_5 <= _T_27720[5];
    conflictPReg_11_6 <= _T_27720[6];
    conflictPReg_11_7 <= _T_27720[7];
    conflictPReg_11_8 <= _T_27720[8];
    conflictPReg_11_9 <= _T_27720[9];
    conflictPReg_11_10 <= _T_27720[10];
    conflictPReg_11_11 <= _T_27720[11];
    conflictPReg_11_12 <= _T_27720[12];
    conflictPReg_11_13 <= _T_27720[13];
    conflictPReg_11_14 <= _T_27720[14];
    conflictPReg_11_15 <= _T_27720[15];
    conflictPReg_12_0 <= _T_28578[0];
    conflictPReg_12_1 <= _T_28578[1];
    conflictPReg_12_2 <= _T_28578[2];
    conflictPReg_12_3 <= _T_28578[3];
    conflictPReg_12_4 <= _T_28578[4];
    conflictPReg_12_5 <= _T_28578[5];
    conflictPReg_12_6 <= _T_28578[6];
    conflictPReg_12_7 <= _T_28578[7];
    conflictPReg_12_8 <= _T_28578[8];
    conflictPReg_12_9 <= _T_28578[9];
    conflictPReg_12_10 <= _T_28578[10];
    conflictPReg_12_11 <= _T_28578[11];
    conflictPReg_12_12 <= _T_28578[12];
    conflictPReg_12_13 <= _T_28578[13];
    conflictPReg_12_14 <= _T_28578[14];
    conflictPReg_12_15 <= _T_28578[15];
    conflictPReg_13_0 <= _T_29436[0];
    conflictPReg_13_1 <= _T_29436[1];
    conflictPReg_13_2 <= _T_29436[2];
    conflictPReg_13_3 <= _T_29436[3];
    conflictPReg_13_4 <= _T_29436[4];
    conflictPReg_13_5 <= _T_29436[5];
    conflictPReg_13_6 <= _T_29436[6];
    conflictPReg_13_7 <= _T_29436[7];
    conflictPReg_13_8 <= _T_29436[8];
    conflictPReg_13_9 <= _T_29436[9];
    conflictPReg_13_10 <= _T_29436[10];
    conflictPReg_13_11 <= _T_29436[11];
    conflictPReg_13_12 <= _T_29436[12];
    conflictPReg_13_13 <= _T_29436[13];
    conflictPReg_13_14 <= _T_29436[14];
    conflictPReg_13_15 <= _T_29436[15];
    conflictPReg_14_0 <= _T_30294[0];
    conflictPReg_14_1 <= _T_30294[1];
    conflictPReg_14_2 <= _T_30294[2];
    conflictPReg_14_3 <= _T_30294[3];
    conflictPReg_14_4 <= _T_30294[4];
    conflictPReg_14_5 <= _T_30294[5];
    conflictPReg_14_6 <= _T_30294[6];
    conflictPReg_14_7 <= _T_30294[7];
    conflictPReg_14_8 <= _T_30294[8];
    conflictPReg_14_9 <= _T_30294[9];
    conflictPReg_14_10 <= _T_30294[10];
    conflictPReg_14_11 <= _T_30294[11];
    conflictPReg_14_12 <= _T_30294[12];
    conflictPReg_14_13 <= _T_30294[13];
    conflictPReg_14_14 <= _T_30294[14];
    conflictPReg_14_15 <= _T_30294[15];
    conflictPReg_15_0 <= _T_31152[0];
    conflictPReg_15_1 <= _T_31152[1];
    conflictPReg_15_2 <= _T_31152[2];
    conflictPReg_15_3 <= _T_31152[3];
    conflictPReg_15_4 <= _T_31152[4];
    conflictPReg_15_5 <= _T_31152[5];
    conflictPReg_15_6 <= _T_31152[6];
    conflictPReg_15_7 <= _T_31152[7];
    conflictPReg_15_8 <= _T_31152[8];
    conflictPReg_15_9 <= _T_31152[9];
    conflictPReg_15_10 <= _T_31152[10];
    conflictPReg_15_11 <= _T_31152[11];
    conflictPReg_15_12 <= _T_31152[12];
    conflictPReg_15_13 <= _T_31152[13];
    conflictPReg_15_14 <= _T_31152[14];
    conflictPReg_15_15 <= _T_31152[15];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_52606[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_52606[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_52606[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_52606[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_52606[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_52606[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_52606[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_52606[7];
    storeAddrNotKnownFlagsPReg_0_8 <= _T_52606[8];
    storeAddrNotKnownFlagsPReg_0_9 <= _T_52606[9];
    storeAddrNotKnownFlagsPReg_0_10 <= _T_52606[10];
    storeAddrNotKnownFlagsPReg_0_11 <= _T_52606[11];
    storeAddrNotKnownFlagsPReg_0_12 <= _T_52606[12];
    storeAddrNotKnownFlagsPReg_0_13 <= _T_52606[13];
    storeAddrNotKnownFlagsPReg_0_14 <= _T_52606[14];
    storeAddrNotKnownFlagsPReg_0_15 <= _T_52606[15];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_53464[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_53464[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_53464[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_53464[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_53464[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_53464[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_53464[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_53464[7];
    storeAddrNotKnownFlagsPReg_1_8 <= _T_53464[8];
    storeAddrNotKnownFlagsPReg_1_9 <= _T_53464[9];
    storeAddrNotKnownFlagsPReg_1_10 <= _T_53464[10];
    storeAddrNotKnownFlagsPReg_1_11 <= _T_53464[11];
    storeAddrNotKnownFlagsPReg_1_12 <= _T_53464[12];
    storeAddrNotKnownFlagsPReg_1_13 <= _T_53464[13];
    storeAddrNotKnownFlagsPReg_1_14 <= _T_53464[14];
    storeAddrNotKnownFlagsPReg_1_15 <= _T_53464[15];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_54322[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_54322[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_54322[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_54322[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_54322[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_54322[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_54322[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_54322[7];
    storeAddrNotKnownFlagsPReg_2_8 <= _T_54322[8];
    storeAddrNotKnownFlagsPReg_2_9 <= _T_54322[9];
    storeAddrNotKnownFlagsPReg_2_10 <= _T_54322[10];
    storeAddrNotKnownFlagsPReg_2_11 <= _T_54322[11];
    storeAddrNotKnownFlagsPReg_2_12 <= _T_54322[12];
    storeAddrNotKnownFlagsPReg_2_13 <= _T_54322[13];
    storeAddrNotKnownFlagsPReg_2_14 <= _T_54322[14];
    storeAddrNotKnownFlagsPReg_2_15 <= _T_54322[15];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_55180[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_55180[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_55180[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_55180[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_55180[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_55180[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_55180[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_55180[7];
    storeAddrNotKnownFlagsPReg_3_8 <= _T_55180[8];
    storeAddrNotKnownFlagsPReg_3_9 <= _T_55180[9];
    storeAddrNotKnownFlagsPReg_3_10 <= _T_55180[10];
    storeAddrNotKnownFlagsPReg_3_11 <= _T_55180[11];
    storeAddrNotKnownFlagsPReg_3_12 <= _T_55180[12];
    storeAddrNotKnownFlagsPReg_3_13 <= _T_55180[13];
    storeAddrNotKnownFlagsPReg_3_14 <= _T_55180[14];
    storeAddrNotKnownFlagsPReg_3_15 <= _T_55180[15];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_56038[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_56038[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_56038[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_56038[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_56038[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_56038[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_56038[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_56038[7];
    storeAddrNotKnownFlagsPReg_4_8 <= _T_56038[8];
    storeAddrNotKnownFlagsPReg_4_9 <= _T_56038[9];
    storeAddrNotKnownFlagsPReg_4_10 <= _T_56038[10];
    storeAddrNotKnownFlagsPReg_4_11 <= _T_56038[11];
    storeAddrNotKnownFlagsPReg_4_12 <= _T_56038[12];
    storeAddrNotKnownFlagsPReg_4_13 <= _T_56038[13];
    storeAddrNotKnownFlagsPReg_4_14 <= _T_56038[14];
    storeAddrNotKnownFlagsPReg_4_15 <= _T_56038[15];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_56896[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_56896[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_56896[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_56896[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_56896[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_56896[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_56896[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_56896[7];
    storeAddrNotKnownFlagsPReg_5_8 <= _T_56896[8];
    storeAddrNotKnownFlagsPReg_5_9 <= _T_56896[9];
    storeAddrNotKnownFlagsPReg_5_10 <= _T_56896[10];
    storeAddrNotKnownFlagsPReg_5_11 <= _T_56896[11];
    storeAddrNotKnownFlagsPReg_5_12 <= _T_56896[12];
    storeAddrNotKnownFlagsPReg_5_13 <= _T_56896[13];
    storeAddrNotKnownFlagsPReg_5_14 <= _T_56896[14];
    storeAddrNotKnownFlagsPReg_5_15 <= _T_56896[15];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_57754[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_57754[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_57754[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_57754[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_57754[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_57754[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_57754[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_57754[7];
    storeAddrNotKnownFlagsPReg_6_8 <= _T_57754[8];
    storeAddrNotKnownFlagsPReg_6_9 <= _T_57754[9];
    storeAddrNotKnownFlagsPReg_6_10 <= _T_57754[10];
    storeAddrNotKnownFlagsPReg_6_11 <= _T_57754[11];
    storeAddrNotKnownFlagsPReg_6_12 <= _T_57754[12];
    storeAddrNotKnownFlagsPReg_6_13 <= _T_57754[13];
    storeAddrNotKnownFlagsPReg_6_14 <= _T_57754[14];
    storeAddrNotKnownFlagsPReg_6_15 <= _T_57754[15];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_58612[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_58612[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_58612[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_58612[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_58612[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_58612[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_58612[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_58612[7];
    storeAddrNotKnownFlagsPReg_7_8 <= _T_58612[8];
    storeAddrNotKnownFlagsPReg_7_9 <= _T_58612[9];
    storeAddrNotKnownFlagsPReg_7_10 <= _T_58612[10];
    storeAddrNotKnownFlagsPReg_7_11 <= _T_58612[11];
    storeAddrNotKnownFlagsPReg_7_12 <= _T_58612[12];
    storeAddrNotKnownFlagsPReg_7_13 <= _T_58612[13];
    storeAddrNotKnownFlagsPReg_7_14 <= _T_58612[14];
    storeAddrNotKnownFlagsPReg_7_15 <= _T_58612[15];
    storeAddrNotKnownFlagsPReg_8_0 <= _T_59470[0];
    storeAddrNotKnownFlagsPReg_8_1 <= _T_59470[1];
    storeAddrNotKnownFlagsPReg_8_2 <= _T_59470[2];
    storeAddrNotKnownFlagsPReg_8_3 <= _T_59470[3];
    storeAddrNotKnownFlagsPReg_8_4 <= _T_59470[4];
    storeAddrNotKnownFlagsPReg_8_5 <= _T_59470[5];
    storeAddrNotKnownFlagsPReg_8_6 <= _T_59470[6];
    storeAddrNotKnownFlagsPReg_8_7 <= _T_59470[7];
    storeAddrNotKnownFlagsPReg_8_8 <= _T_59470[8];
    storeAddrNotKnownFlagsPReg_8_9 <= _T_59470[9];
    storeAddrNotKnownFlagsPReg_8_10 <= _T_59470[10];
    storeAddrNotKnownFlagsPReg_8_11 <= _T_59470[11];
    storeAddrNotKnownFlagsPReg_8_12 <= _T_59470[12];
    storeAddrNotKnownFlagsPReg_8_13 <= _T_59470[13];
    storeAddrNotKnownFlagsPReg_8_14 <= _T_59470[14];
    storeAddrNotKnownFlagsPReg_8_15 <= _T_59470[15];
    storeAddrNotKnownFlagsPReg_9_0 <= _T_60328[0];
    storeAddrNotKnownFlagsPReg_9_1 <= _T_60328[1];
    storeAddrNotKnownFlagsPReg_9_2 <= _T_60328[2];
    storeAddrNotKnownFlagsPReg_9_3 <= _T_60328[3];
    storeAddrNotKnownFlagsPReg_9_4 <= _T_60328[4];
    storeAddrNotKnownFlagsPReg_9_5 <= _T_60328[5];
    storeAddrNotKnownFlagsPReg_9_6 <= _T_60328[6];
    storeAddrNotKnownFlagsPReg_9_7 <= _T_60328[7];
    storeAddrNotKnownFlagsPReg_9_8 <= _T_60328[8];
    storeAddrNotKnownFlagsPReg_9_9 <= _T_60328[9];
    storeAddrNotKnownFlagsPReg_9_10 <= _T_60328[10];
    storeAddrNotKnownFlagsPReg_9_11 <= _T_60328[11];
    storeAddrNotKnownFlagsPReg_9_12 <= _T_60328[12];
    storeAddrNotKnownFlagsPReg_9_13 <= _T_60328[13];
    storeAddrNotKnownFlagsPReg_9_14 <= _T_60328[14];
    storeAddrNotKnownFlagsPReg_9_15 <= _T_60328[15];
    storeAddrNotKnownFlagsPReg_10_0 <= _T_61186[0];
    storeAddrNotKnownFlagsPReg_10_1 <= _T_61186[1];
    storeAddrNotKnownFlagsPReg_10_2 <= _T_61186[2];
    storeAddrNotKnownFlagsPReg_10_3 <= _T_61186[3];
    storeAddrNotKnownFlagsPReg_10_4 <= _T_61186[4];
    storeAddrNotKnownFlagsPReg_10_5 <= _T_61186[5];
    storeAddrNotKnownFlagsPReg_10_6 <= _T_61186[6];
    storeAddrNotKnownFlagsPReg_10_7 <= _T_61186[7];
    storeAddrNotKnownFlagsPReg_10_8 <= _T_61186[8];
    storeAddrNotKnownFlagsPReg_10_9 <= _T_61186[9];
    storeAddrNotKnownFlagsPReg_10_10 <= _T_61186[10];
    storeAddrNotKnownFlagsPReg_10_11 <= _T_61186[11];
    storeAddrNotKnownFlagsPReg_10_12 <= _T_61186[12];
    storeAddrNotKnownFlagsPReg_10_13 <= _T_61186[13];
    storeAddrNotKnownFlagsPReg_10_14 <= _T_61186[14];
    storeAddrNotKnownFlagsPReg_10_15 <= _T_61186[15];
    storeAddrNotKnownFlagsPReg_11_0 <= _T_62044[0];
    storeAddrNotKnownFlagsPReg_11_1 <= _T_62044[1];
    storeAddrNotKnownFlagsPReg_11_2 <= _T_62044[2];
    storeAddrNotKnownFlagsPReg_11_3 <= _T_62044[3];
    storeAddrNotKnownFlagsPReg_11_4 <= _T_62044[4];
    storeAddrNotKnownFlagsPReg_11_5 <= _T_62044[5];
    storeAddrNotKnownFlagsPReg_11_6 <= _T_62044[6];
    storeAddrNotKnownFlagsPReg_11_7 <= _T_62044[7];
    storeAddrNotKnownFlagsPReg_11_8 <= _T_62044[8];
    storeAddrNotKnownFlagsPReg_11_9 <= _T_62044[9];
    storeAddrNotKnownFlagsPReg_11_10 <= _T_62044[10];
    storeAddrNotKnownFlagsPReg_11_11 <= _T_62044[11];
    storeAddrNotKnownFlagsPReg_11_12 <= _T_62044[12];
    storeAddrNotKnownFlagsPReg_11_13 <= _T_62044[13];
    storeAddrNotKnownFlagsPReg_11_14 <= _T_62044[14];
    storeAddrNotKnownFlagsPReg_11_15 <= _T_62044[15];
    storeAddrNotKnownFlagsPReg_12_0 <= _T_62902[0];
    storeAddrNotKnownFlagsPReg_12_1 <= _T_62902[1];
    storeAddrNotKnownFlagsPReg_12_2 <= _T_62902[2];
    storeAddrNotKnownFlagsPReg_12_3 <= _T_62902[3];
    storeAddrNotKnownFlagsPReg_12_4 <= _T_62902[4];
    storeAddrNotKnownFlagsPReg_12_5 <= _T_62902[5];
    storeAddrNotKnownFlagsPReg_12_6 <= _T_62902[6];
    storeAddrNotKnownFlagsPReg_12_7 <= _T_62902[7];
    storeAddrNotKnownFlagsPReg_12_8 <= _T_62902[8];
    storeAddrNotKnownFlagsPReg_12_9 <= _T_62902[9];
    storeAddrNotKnownFlagsPReg_12_10 <= _T_62902[10];
    storeAddrNotKnownFlagsPReg_12_11 <= _T_62902[11];
    storeAddrNotKnownFlagsPReg_12_12 <= _T_62902[12];
    storeAddrNotKnownFlagsPReg_12_13 <= _T_62902[13];
    storeAddrNotKnownFlagsPReg_12_14 <= _T_62902[14];
    storeAddrNotKnownFlagsPReg_12_15 <= _T_62902[15];
    storeAddrNotKnownFlagsPReg_13_0 <= _T_63760[0];
    storeAddrNotKnownFlagsPReg_13_1 <= _T_63760[1];
    storeAddrNotKnownFlagsPReg_13_2 <= _T_63760[2];
    storeAddrNotKnownFlagsPReg_13_3 <= _T_63760[3];
    storeAddrNotKnownFlagsPReg_13_4 <= _T_63760[4];
    storeAddrNotKnownFlagsPReg_13_5 <= _T_63760[5];
    storeAddrNotKnownFlagsPReg_13_6 <= _T_63760[6];
    storeAddrNotKnownFlagsPReg_13_7 <= _T_63760[7];
    storeAddrNotKnownFlagsPReg_13_8 <= _T_63760[8];
    storeAddrNotKnownFlagsPReg_13_9 <= _T_63760[9];
    storeAddrNotKnownFlagsPReg_13_10 <= _T_63760[10];
    storeAddrNotKnownFlagsPReg_13_11 <= _T_63760[11];
    storeAddrNotKnownFlagsPReg_13_12 <= _T_63760[12];
    storeAddrNotKnownFlagsPReg_13_13 <= _T_63760[13];
    storeAddrNotKnownFlagsPReg_13_14 <= _T_63760[14];
    storeAddrNotKnownFlagsPReg_13_15 <= _T_63760[15];
    storeAddrNotKnownFlagsPReg_14_0 <= _T_64618[0];
    storeAddrNotKnownFlagsPReg_14_1 <= _T_64618[1];
    storeAddrNotKnownFlagsPReg_14_2 <= _T_64618[2];
    storeAddrNotKnownFlagsPReg_14_3 <= _T_64618[3];
    storeAddrNotKnownFlagsPReg_14_4 <= _T_64618[4];
    storeAddrNotKnownFlagsPReg_14_5 <= _T_64618[5];
    storeAddrNotKnownFlagsPReg_14_6 <= _T_64618[6];
    storeAddrNotKnownFlagsPReg_14_7 <= _T_64618[7];
    storeAddrNotKnownFlagsPReg_14_8 <= _T_64618[8];
    storeAddrNotKnownFlagsPReg_14_9 <= _T_64618[9];
    storeAddrNotKnownFlagsPReg_14_10 <= _T_64618[10];
    storeAddrNotKnownFlagsPReg_14_11 <= _T_64618[11];
    storeAddrNotKnownFlagsPReg_14_12 <= _T_64618[12];
    storeAddrNotKnownFlagsPReg_14_13 <= _T_64618[13];
    storeAddrNotKnownFlagsPReg_14_14 <= _T_64618[14];
    storeAddrNotKnownFlagsPReg_14_15 <= _T_64618[15];
    storeAddrNotKnownFlagsPReg_15_0 <= _T_65476[0];
    storeAddrNotKnownFlagsPReg_15_1 <= _T_65476[1];
    storeAddrNotKnownFlagsPReg_15_2 <= _T_65476[2];
    storeAddrNotKnownFlagsPReg_15_3 <= _T_65476[3];
    storeAddrNotKnownFlagsPReg_15_4 <= _T_65476[4];
    storeAddrNotKnownFlagsPReg_15_5 <= _T_65476[5];
    storeAddrNotKnownFlagsPReg_15_6 <= _T_65476[6];
    storeAddrNotKnownFlagsPReg_15_7 <= _T_65476[7];
    storeAddrNotKnownFlagsPReg_15_8 <= _T_65476[8];
    storeAddrNotKnownFlagsPReg_15_9 <= _T_65476[9];
    storeAddrNotKnownFlagsPReg_15_10 <= _T_65476[10];
    storeAddrNotKnownFlagsPReg_15_11 <= _T_65476[11];
    storeAddrNotKnownFlagsPReg_15_12 <= _T_65476[12];
    storeAddrNotKnownFlagsPReg_15_13 <= _T_65476[13];
    storeAddrNotKnownFlagsPReg_15_14 <= _T_65476[14];
    storeAddrNotKnownFlagsPReg_15_15 <= _T_65476[15];
    shiftedStoreDataKnownPReg_0 <= _T_5972[0];
    shiftedStoreDataKnownPReg_1 <= _T_5972[1];
    shiftedStoreDataKnownPReg_2 <= _T_5972[2];
    shiftedStoreDataKnownPReg_3 <= _T_5972[3];
    shiftedStoreDataKnownPReg_4 <= _T_5972[4];
    shiftedStoreDataKnownPReg_5 <= _T_5972[5];
    shiftedStoreDataKnownPReg_6 <= _T_5972[6];
    shiftedStoreDataKnownPReg_7 <= _T_5972[7];
    shiftedStoreDataKnownPReg_8 <= _T_5972[8];
    shiftedStoreDataKnownPReg_9 <= _T_5972[9];
    shiftedStoreDataKnownPReg_10 <= _T_5972[10];
    shiftedStoreDataKnownPReg_11 <= _T_5972[11];
    shiftedStoreDataKnownPReg_12 <= _T_5972[12];
    shiftedStoreDataKnownPReg_13 <= _T_5972[13];
    shiftedStoreDataKnownPReg_14 <= _T_5972[14];
    shiftedStoreDataKnownPReg_15 <= _T_5972[15];
    shiftedStoreDataQPreg_0 <= _T_5115[31:0];
    shiftedStoreDataQPreg_1 <= _T_5115[63:32];
    shiftedStoreDataQPreg_2 <= _T_5115[95:64];
    shiftedStoreDataQPreg_3 <= _T_5115[127:96];
    shiftedStoreDataQPreg_4 <= _T_5115[159:128];
    shiftedStoreDataQPreg_5 <= _T_5115[191:160];
    shiftedStoreDataQPreg_6 <= _T_5115[223:192];
    shiftedStoreDataQPreg_7 <= _T_5115[255:224];
    shiftedStoreDataQPreg_8 <= _T_5115[287:256];
    shiftedStoreDataQPreg_9 <= _T_5115[319:288];
    shiftedStoreDataQPreg_10 <= _T_5115[351:320];
    shiftedStoreDataQPreg_11 <= _T_5115[383:352];
    shiftedStoreDataQPreg_12 <= _T_5115[415:384];
    shiftedStoreDataQPreg_13 <= _T_5115[447:416];
    shiftedStoreDataQPreg_14 <= _T_5115[479:448];
    shiftedStoreDataQPreg_15 <= _T_5115[511:480];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    addrKnownPReg_8 <= addrKnown_8;
    addrKnownPReg_9 <= addrKnown_9;
    addrKnownPReg_10 <= addrKnown_10;
    addrKnownPReg_11 <= addrKnown_11;
    addrKnownPReg_12 <= addrKnown_12;
    addrKnownPReg_13 <= addrKnown_13;
    addrKnownPReg_14 <= addrKnown_14;
    addrKnownPReg_15 <= addrKnown_15;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    dataKnownPReg_8 <= dataKnown_8;
    dataKnownPReg_9 <= dataKnown_9;
    dataKnownPReg_10 <= dataKnown_10;
    dataKnownPReg_11 <= dataKnown_11;
    dataKnownPReg_12 <= dataKnown_12;
    dataKnownPReg_13 <= dataKnown_13;
    dataKnownPReg_14 <= dataKnown_14;
    dataKnownPReg_15 <= dataKnown_15;
    if (reset) begin
      prevPriorityRequest_15 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_15 <= priorityLoadRequest_15;
      end else begin
        prevPriorityRequest_15 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_14 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_14 <= priorityLoadRequest_14;
      end else begin
        prevPriorityRequest_14 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_13 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_13 <= priorityLoadRequest_13;
      end else begin
        prevPriorityRequest_13 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_12 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_12 <= priorityLoadRequest_12;
      end else begin
        prevPriorityRequest_12 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_11 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_11 <= priorityLoadRequest_11;
      end else begin
        prevPriorityRequest_11 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_10 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_10 <= priorityLoadRequest_10;
      end else begin
        prevPriorityRequest_10 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_9 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_9 <= priorityLoadRequest_9;
      end else begin
        prevPriorityRequest_9 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_8 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_8 <= priorityLoadRequest_8;
      end else begin
        prevPriorityRequest_8 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_7 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_7 <= priorityLoadRequest_7;
      end else begin
        prevPriorityRequest_7 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_6 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_6 <= priorityLoadRequest_6;
      end else begin
        prevPriorityRequest_6 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_5 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_5 <= priorityLoadRequest_5;
      end else begin
        prevPriorityRequest_5 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_4 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_4 <= priorityLoadRequest_4;
      end else begin
        prevPriorityRequest_4 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_3 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_3 <= priorityLoadRequest_3;
      end else begin
        prevPriorityRequest_3 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_2 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_2 <= priorityLoadRequest_2;
      end else begin
        prevPriorityRequest_2 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_1 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_1 <= priorityLoadRequest_1;
      end else begin
        prevPriorityRequest_1 <= 1'h0;
      end
    end
    if (reset) begin
      prevPriorityRequest_0 <= 1'h0;
    end else begin
      if (io_memIsReadyForLoads) begin
        prevPriorityRequest_0 <= priorityLoadRequest_0;
      end else begin
        prevPriorityRequest_0 <= 1'h0;
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_A( // @[:@42439.2]
  output [3:0] io_bbLoadOffsets_0, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_1, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_2, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_3, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_4, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_5, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_6, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_7, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_8, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_9, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_10, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_11, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_12, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_13, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_14, // @[:@42442.4]
  output [3:0] io_bbLoadOffsets_15, // @[:@42442.4]
  output       io_bbNumLoads, // @[:@42442.4]
  input  [3:0] io_loadTail, // @[:@42442.4]
  input  [3:0] io_loadHead, // @[:@42442.4]
  input        io_loadEmpty, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_0, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_1, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_2, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_3, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_4, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_5, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_6, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_7, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_8, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_9, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_10, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_11, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_12, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_13, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_14, // @[:@42442.4]
  output [3:0] io_bbStoreOffsets_15, // @[:@42442.4]
  output       io_bbNumStores, // @[:@42442.4]
  input  [3:0] io_storeTail, // @[:@42442.4]
  input  [3:0] io_storeHead, // @[:@42442.4]
  input        io_storeEmpty, // @[:@42442.4]
  output       io_bbStart, // @[:@42442.4]
  input        io_bbStartSignals_0, // @[:@42442.4]
  input        io_bbStartSignals_1, // @[:@42442.4]
  output       io_readyToPrevious_0, // @[:@42442.4]
  output       io_readyToPrevious_1, // @[:@42442.4]
  output       io_loadPortsEnable_0, // @[:@42442.4]
  output       io_storePortsEnable_0 // @[:@42442.4]
);
  wire  _T_244; // @[GroupAllocator.scala 42:25:@42445.4]
  wire  _T_245; // @[GroupAllocator.scala 42:16:@42446.4]
  wire [4:0] _GEN_68; // @[GroupAllocator.scala 43:36:@42448.6]
  wire [5:0] _T_247; // @[GroupAllocator.scala 43:36:@42448.6]
  wire [5:0] _T_248; // @[GroupAllocator.scala 43:36:@42449.6]
  wire [4:0] _T_249; // @[GroupAllocator.scala 43:36:@42450.6]
  wire [4:0] _GEN_69; // @[GroupAllocator.scala 43:43:@42451.6]
  wire [5:0] _T_250; // @[GroupAllocator.scala 43:43:@42451.6]
  wire [4:0] _T_251; // @[GroupAllocator.scala 43:43:@42452.6]
  wire [4:0] _T_252; // @[GroupAllocator.scala 45:22:@42456.6]
  wire [4:0] _T_253; // @[GroupAllocator.scala 45:22:@42457.6]
  wire [3:0] _T_254; // @[GroupAllocator.scala 45:22:@42458.6]
  wire [4:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@42447.4]
  wire  _T_256; // @[GroupAllocator.scala 42:25:@42462.4]
  wire  _T_257; // @[GroupAllocator.scala 42:16:@42463.4]
  wire [4:0] _GEN_70; // @[GroupAllocator.scala 43:36:@42465.6]
  wire [5:0] _T_259; // @[GroupAllocator.scala 43:36:@42465.6]
  wire [5:0] _T_260; // @[GroupAllocator.scala 43:36:@42466.6]
  wire [4:0] _T_261; // @[GroupAllocator.scala 43:36:@42467.6]
  wire [4:0] _GEN_71; // @[GroupAllocator.scala 43:43:@42468.6]
  wire [5:0] _T_262; // @[GroupAllocator.scala 43:43:@42468.6]
  wire [4:0] _T_263; // @[GroupAllocator.scala 43:43:@42469.6]
  wire [4:0] _T_264; // @[GroupAllocator.scala 45:22:@42473.6]
  wire [4:0] _T_265; // @[GroupAllocator.scala 45:22:@42474.6]
  wire [3:0] _T_266; // @[GroupAllocator.scala 45:22:@42475.6]
  wire [4:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@42464.4]
  wire  possibleAllocations_0; // @[GroupAllocator.scala 56:106:@42489.4]
  wire  possibleAllocations_1; // @[GroupAllocator.scala 56:106:@42490.4]
  wire  allocatedBBIdx; // @[Mux.scala 31:69:@42494.4]
  wire  _T_300; // @[GroupAllocator.scala 69:43:@42498.4]
  wire  _T_476; // @[Mux.scala 46:16:@42647.6]
  wire [5:0] _T_898; // @[GroupAllocator.scala 110:34:@42808.6]
  wire [4:0] _T_899; // @[GroupAllocator.scala 110:34:@42809.6]
  wire [5:0] _T_901; // @[GroupAllocator.scala 110:55:@42810.6]
  wire [5:0] _T_902; // @[GroupAllocator.scala 110:55:@42811.6]
  wire [4:0] _T_903; // @[GroupAllocator.scala 110:55:@42812.6]
  wire [5:0] _T_905; // @[util.scala 10:8:@42813.6]
  wire [5:0] _GEN_0; // @[util.scala 10:14:@42814.6]
  wire [4:0] _T_906; // @[util.scala 10:14:@42814.6]
  wire [3:0] _T_1156; // @[GroupAllocator.scala 110:90:@42976.6 GroupAllocator.scala 110:90:@42977.6]
  wire [3:0] _T_1390_0; // @[Mux.scala 46:16:@43131.6]
  wire [3:0] _T_1427_0; // @[Mux.scala 46:16:@43133.6]
  wire [5:0] _T_1504; // @[GroupAllocator.scala 115:33:@43167.6]
  wire [4:0] _T_1505; // @[GroupAllocator.scala 115:33:@43168.6]
  wire [5:0] _T_1507; // @[GroupAllocator.scala 115:54:@43169.6]
  wire [5:0] _T_1508; // @[GroupAllocator.scala 115:54:@43170.6]
  wire [4:0] _T_1509; // @[GroupAllocator.scala 115:54:@43171.6]
  wire [5:0] _T_1511; // @[util.scala 10:8:@43172.6]
  wire [5:0] _GEN_1; // @[util.scala 10:14:@43173.6]
  wire [4:0] _T_1512; // @[util.scala 10:14:@43173.6]
  wire [3:0] _T_1762; // @[GroupAllocator.scala 115:89:@43335.6 GroupAllocator.scala 115:89:@43336.6]
  wire [3:0] _T_1996_0; // @[Mux.scala 46:16:@43490.6]
  wire [3:0] _T_2033_0; // @[Mux.scala 46:16:@43492.6]
  assign _T_244 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@42445.4]
  assign _T_245 = io_loadEmpty | _T_244; // @[GroupAllocator.scala 42:16:@42446.4]
  assign _GEN_68 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@42448.6]
  assign _T_247 = 5'h10 - _GEN_68; // @[GroupAllocator.scala 43:36:@42448.6]
  assign _T_248 = $unsigned(_T_247); // @[GroupAllocator.scala 43:36:@42449.6]
  assign _T_249 = _T_248[4:0]; // @[GroupAllocator.scala 43:36:@42450.6]
  assign _GEN_69 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@42451.6]
  assign _T_250 = _T_249 + _GEN_69; // @[GroupAllocator.scala 43:43:@42451.6]
  assign _T_251 = _T_249 + _GEN_69; // @[GroupAllocator.scala 43:43:@42452.6]
  assign _T_252 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@42456.6]
  assign _T_253 = $unsigned(_T_252); // @[GroupAllocator.scala 45:22:@42457.6]
  assign _T_254 = _T_253[3:0]; // @[GroupAllocator.scala 45:22:@42458.6]
  assign emptyLoadSlots = _T_245 ? _T_251 : {{1'd0}, _T_254}; // @[GroupAllocator.scala 42:34:@42447.4]
  assign _T_256 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@42462.4]
  assign _T_257 = io_storeEmpty | _T_256; // @[GroupAllocator.scala 42:16:@42463.4]
  assign _GEN_70 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@42465.6]
  assign _T_259 = 5'h10 - _GEN_70; // @[GroupAllocator.scala 43:36:@42465.6]
  assign _T_260 = $unsigned(_T_259); // @[GroupAllocator.scala 43:36:@42466.6]
  assign _T_261 = _T_260[4:0]; // @[GroupAllocator.scala 43:36:@42467.6]
  assign _GEN_71 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@42468.6]
  assign _T_262 = _T_261 + _GEN_71; // @[GroupAllocator.scala 43:43:@42468.6]
  assign _T_263 = _T_261 + _GEN_71; // @[GroupAllocator.scala 43:43:@42469.6]
  assign _T_264 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@42473.6]
  assign _T_265 = $unsigned(_T_264); // @[GroupAllocator.scala 45:22:@42474.6]
  assign _T_266 = _T_265[3:0]; // @[GroupAllocator.scala 45:22:@42475.6]
  assign emptyStoreSlots = _T_257 ? _T_263 : {{1'd0}, _T_266}; // @[GroupAllocator.scala 42:34:@42464.4]
  assign possibleAllocations_0 = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 56:106:@42489.4]
  assign possibleAllocations_1 = io_readyToPrevious_1 & io_bbStartSignals_1; // @[GroupAllocator.scala 56:106:@42490.4]
  assign allocatedBBIdx = possibleAllocations_0 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@42494.4]
  assign _T_300 = 1'h0 == allocatedBBIdx; // @[GroupAllocator.scala 69:43:@42498.4]
  assign _T_476 = _T_300 ? 1'h0 : allocatedBBIdx; // @[Mux.scala 46:16:@42647.6]
  assign _T_898 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@42808.6]
  assign _T_899 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@42809.6]
  assign _T_901 = _T_899 - 5'h1; // @[GroupAllocator.scala 110:55:@42810.6]
  assign _T_902 = $unsigned(_T_901); // @[GroupAllocator.scala 110:55:@42811.6]
  assign _T_903 = _T_902[4:0]; // @[GroupAllocator.scala 110:55:@42812.6]
  assign _T_905 = {{1'd0}, _T_903}; // @[util.scala 10:8:@42813.6]
  assign _GEN_0 = _T_905 % 6'h10; // @[util.scala 10:14:@42814.6]
  assign _T_906 = _GEN_0[4:0]; // @[util.scala 10:14:@42814.6]
  assign _T_1156 = _T_906[3:0]; // @[GroupAllocator.scala 110:90:@42976.6 GroupAllocator.scala 110:90:@42977.6]
  assign _T_1390_0 = allocatedBBIdx ? _T_1156 : 4'h0; // @[Mux.scala 46:16:@43131.6]
  assign _T_1427_0 = _T_300 ? _T_1156 : _T_1390_0; // @[Mux.scala 46:16:@43133.6]
  assign _T_1504 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@43167.6]
  assign _T_1505 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@43168.6]
  assign _T_1507 = _T_1505 - 5'h1; // @[GroupAllocator.scala 115:54:@43169.6]
  assign _T_1508 = $unsigned(_T_1507); // @[GroupAllocator.scala 115:54:@43170.6]
  assign _T_1509 = _T_1508[4:0]; // @[GroupAllocator.scala 115:54:@43171.6]
  assign _T_1511 = {{1'd0}, _T_1509}; // @[util.scala 10:8:@43172.6]
  assign _GEN_1 = _T_1511 % 6'h10; // @[util.scala 10:14:@43173.6]
  assign _T_1512 = _GEN_1[4:0]; // @[util.scala 10:14:@43173.6]
  assign _T_1762 = _T_1512[3:0]; // @[GroupAllocator.scala 115:89:@43335.6 GroupAllocator.scala 115:89:@43336.6]
  assign _T_1996_0 = allocatedBBIdx ? _T_1762 : 4'h0; // @[Mux.scala 46:16:@43490.6]
  assign _T_2033_0 = _T_300 ? _T_1762 : _T_1996_0; // @[Mux.scala 46:16:@43492.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42589.4 GroupAllocator.scala 106:22:@43134.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42590.4 GroupAllocator.scala 106:22:@43135.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42591.4 GroupAllocator.scala 106:22:@43136.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42592.4 GroupAllocator.scala 106:22:@43137.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42593.4 GroupAllocator.scala 106:22:@43138.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42594.4 GroupAllocator.scala 106:22:@43139.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42595.4 GroupAllocator.scala 106:22:@43140.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42596.4 GroupAllocator.scala 106:22:@43141.6]
  assign io_bbLoadOffsets_8 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42597.4 GroupAllocator.scala 106:22:@43142.6]
  assign io_bbLoadOffsets_9 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42598.4 GroupAllocator.scala 106:22:@43143.6]
  assign io_bbLoadOffsets_10 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42599.4 GroupAllocator.scala 106:22:@43144.6]
  assign io_bbLoadOffsets_11 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42600.4 GroupAllocator.scala 106:22:@43145.6]
  assign io_bbLoadOffsets_12 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42601.4 GroupAllocator.scala 106:22:@43146.6]
  assign io_bbLoadOffsets_13 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42602.4 GroupAllocator.scala 106:22:@43147.6]
  assign io_bbLoadOffsets_14 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42603.4 GroupAllocator.scala 106:22:@43148.6]
  assign io_bbLoadOffsets_15 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42604.4 GroupAllocator.scala 106:22:@43149.6]
  assign io_bbNumLoads = io_bbStart ? _T_300 : 1'h0; // @[GroupAllocator.scala 85:17:@42504.4 GroupAllocator.scala 93:19:@42643.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42622.4 GroupAllocator.scala 111:23:@43493.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42623.4 GroupAllocator.scala 111:23:@43494.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42624.4 GroupAllocator.scala 111:23:@43495.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42625.4 GroupAllocator.scala 111:23:@43496.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42626.4 GroupAllocator.scala 111:23:@43497.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42627.4 GroupAllocator.scala 111:23:@43498.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42628.4 GroupAllocator.scala 111:23:@43499.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42629.4 GroupAllocator.scala 111:23:@43500.6]
  assign io_bbStoreOffsets_8 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42630.4 GroupAllocator.scala 111:23:@43501.6]
  assign io_bbStoreOffsets_9 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42631.4 GroupAllocator.scala 111:23:@43502.6]
  assign io_bbStoreOffsets_10 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42632.4 GroupAllocator.scala 111:23:@43503.6]
  assign io_bbStoreOffsets_11 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42633.4 GroupAllocator.scala 111:23:@43504.6]
  assign io_bbStoreOffsets_12 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42634.4 GroupAllocator.scala 111:23:@43505.6]
  assign io_bbStoreOffsets_13 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42635.4 GroupAllocator.scala 111:23:@43506.6]
  assign io_bbStoreOffsets_14 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42636.4 GroupAllocator.scala 111:23:@43507.6]
  assign io_bbStoreOffsets_15 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42637.4 GroupAllocator.scala 111:23:@43508.6]
  assign io_bbNumStores = io_bbStart ? _T_476 : 1'h0; // @[GroupAllocator.scala 86:18:@42505.4 GroupAllocator.scala 94:20:@42648.6]
  assign io_bbStart = possibleAllocations_0 | possibleAllocations_1; // @[GroupAllocator.scala 59:14:@42497.4]
  assign io_readyToPrevious_0 = 5'h1 <= emptyLoadSlots; // @[GroupAllocator.scala 53:22:@42487.4]
  assign io_readyToPrevious_1 = 5'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 53:22:@42488.4]
  assign io_loadPortsEnable_0 = _T_300 & io_bbStart; // @[GroupAllocator.scala 69:29:@42500.4]
  assign io_storePortsEnable_0 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 78:30:@42503.4]
endmodule
module LOAD_PORT_LSQ_A( // @[:@43511.2]
  input         clock, // @[:@43512.4]
  input         reset, // @[:@43513.4]
  output        io_addrFromPrev_ready, // @[:@43514.4]
  input         io_addrFromPrev_valid, // @[:@43514.4]
  input  [31:0] io_addrFromPrev_bits, // @[:@43514.4]
  input         io_portEnable, // @[:@43514.4]
  input         io_dataToNext_ready, // @[:@43514.4]
  output        io_dataToNext_valid, // @[:@43514.4]
  output [31:0] io_dataToNext_bits, // @[:@43514.4]
  output        io_loadAddrEnable, // @[:@43514.4]
  output [31:0] io_addrToLoadQueue, // @[:@43514.4]
  output        io_dataFromLoadQueue_ready, // @[:@43514.4]
  input         io_dataFromLoadQueue_valid, // @[:@43514.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@43514.4]
);
  reg [4:0] cnt; // @[LoadPort.scala 23:20:@43516.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@43517.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@43518.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@43519.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@43520.4]
  wire [5:0] _T_50; // @[LoadPort.scala 27:16:@43522.6]
  wire [4:0] _T_51; // @[LoadPort.scala 27:16:@43523.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@43527.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@43528.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@43529.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@43530.6]
  wire [5:0] _T_59; // @[LoadPort.scala 29:16:@43532.8]
  wire [5:0] _T_60; // @[LoadPort.scala 29:16:@43533.8]
  wire [4:0] _T_61; // @[LoadPort.scala 29:16:@43534.8]
  wire [4:0] _GEN_0; // @[LoadPort.scala 28:66:@43531.6]
  wire [4:0] _GEN_1; // @[LoadPort.scala 26:75:@43521.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@43538.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@43517.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@43518.4]
  assign _T_47 = cnt != 5'h10; // @[LoadPort.scala 26:51:@43519.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@43520.4]
  assign _T_50 = cnt + 5'h1; // @[LoadPort.scala 27:16:@43522.6]
  assign _T_51 = cnt + 5'h1; // @[LoadPort.scala 27:16:@43523.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@43527.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@43528.6]
  assign _T_56 = cnt != 5'h0; // @[LoadPort.scala 28:57:@43529.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@43530.6]
  assign _T_59 = cnt - 5'h1; // @[LoadPort.scala 29:16:@43532.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@43533.8]
  assign _T_61 = _T_60[4:0]; // @[LoadPort.scala 29:16:@43534.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@43531.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@43521.4]
  assign _T_63 = cnt > 5'h0; // @[LoadPort.scala 33:28:@43538.4]
  assign io_addrFromPrev_ready = cnt > 5'h0; // @[LoadPort.scala 34:25:@43542.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@43544.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@43543.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@43540.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@43537.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@43545.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_A( // @[:@43547.2]
  input         clock, // @[:@43548.4]
  input         reset, // @[:@43549.4]
  output        io_dataFromPrev_ready, // @[:@43550.4]
  input         io_dataFromPrev_valid, // @[:@43550.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@43550.4]
  input         io_portEnable, // @[:@43550.4]
  output        io_storeDataEnable, // @[:@43550.4]
  output [31:0] io_dataToStoreQueue // @[:@43550.4]
);
  reg [4:0] cnt; // @[StoreDataPort.scala 21:20:@43552.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@43553.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@43554.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@43555.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@43556.4]
  wire [5:0] _T_32; // @[StoreDataPort.scala 25:16:@43558.6]
  wire [4:0] _T_33; // @[StoreDataPort.scala 25:16:@43559.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@43563.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@43564.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@43565.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@43566.6]
  wire [5:0] _T_41; // @[StoreDataPort.scala 27:16:@43568.8]
  wire [5:0] _T_42; // @[StoreDataPort.scala 27:16:@43569.8]
  wire [4:0] _T_43; // @[StoreDataPort.scala 27:16:@43570.8]
  wire [4:0] _GEN_0; // @[StoreDataPort.scala 26:67:@43567.6]
  wire [4:0] _GEN_1; // @[StoreDataPort.scala 24:76:@43557.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@43574.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@43553.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@43554.4]
  assign _T_29 = cnt != 5'h10; // @[StoreDataPort.scala 24:52:@43555.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@43556.4]
  assign _T_32 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@43558.6]
  assign _T_33 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@43559.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@43563.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@43564.6]
  assign _T_38 = cnt != 5'h0; // @[StoreDataPort.scala 26:58:@43565.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@43566.6]
  assign _T_41 = cnt - 5'h1; // @[StoreDataPort.scala 27:16:@43568.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@43569.8]
  assign _T_43 = _T_42[4:0]; // @[StoreDataPort.scala 27:16:@43570.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@43567.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@43557.4]
  assign _T_45 = cnt > 5'h0; // @[StoreDataPort.scala 31:29:@43574.4]
  assign io_dataFromPrev_ready = cnt > 5'h0; // @[StoreDataPort.scala 32:25:@43578.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@43576.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@43573.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_A( // @[:@43613.2]
  input         clock, // @[:@43614.4]
  input         reset, // @[:@43615.4]
  output [31:0] io_storeDataOut, // @[:@43616.4]
  output [31:0] io_storeAddrOut, // @[:@43616.4]
  output        io_storeEnable, // @[:@43616.4]
  input         io_memIsReadyForStores, // @[:@43616.4]
  input  [31:0] io_loadDataIn, // @[:@43616.4]
  output [31:0] io_loadAddrOut, // @[:@43616.4]
  output        io_loadEnable, // @[:@43616.4]
  input         io_memIsReadyForLoads, // @[:@43616.4]
  input         io_bbpValids_0, // @[:@43616.4]
  input         io_bbpValids_1, // @[:@43616.4]
  output        io_bbReadyToPrevs_0, // @[:@43616.4]
  output        io_bbReadyToPrevs_1, // @[:@43616.4]
  output        io_rdPortsPrev_0_ready, // @[:@43616.4]
  input         io_rdPortsPrev_0_valid, // @[:@43616.4]
  input  [31:0] io_rdPortsPrev_0_bits, // @[:@43616.4]
  input         io_rdPortsNext_0_ready, // @[:@43616.4]
  output        io_rdPortsNext_0_valid, // @[:@43616.4]
  output [31:0] io_rdPortsNext_0_bits, // @[:@43616.4]
  output        io_wrAddrPorts_0_ready, // @[:@43616.4]
  input         io_wrAddrPorts_0_valid, // @[:@43616.4]
  input  [31:0] io_wrAddrPorts_0_bits, // @[:@43616.4]
  output        io_wrDataPorts_0_ready, // @[:@43616.4]
  input         io_wrDataPorts_0_valid, // @[:@43616.4]
  input  [31:0] io_wrDataPorts_0_bits, // @[:@43616.4]
  output        io_Empty_Valid // @[:@43616.4]
);
  wire  storeQ_clock; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_reset; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_bbStart; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_bbStoreOffsets_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_bbNumStores; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_storeTail; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_storeHead; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeEmpty; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_loadTail; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [3:0] storeQ_io_loadHead; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadEmpty; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadAddressDone_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_loadDataDone_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_loadAddressQueue_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_addressFromStorePorts_0; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 72:22:@43647.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  storeQ_io_memIsReadyForStores; // @[LSQBRAM.scala 72:22:@43647.4]
  wire  loadQ_clock; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_reset; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_bbStart; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_bbLoadOffsets_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_bbNumLoads; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_loadTail; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_loadHead; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadEmpty; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_storeTail; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] loadQ_io_storeHead; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeEmpty; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeAddrDone_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_storeDataDone_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_storeDataQueue_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_addrFromLoadPorts_0; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [31:0] loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 73:21:@43650.4]
  wire  loadQ_io_memIsReadyForLoads; // @[LSQBRAM.scala 73:21:@43650.4]
  wire [3:0] GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_bbNumLoads; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_loadTail; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_loadHead; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_loadEmpty; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_bbNumStores; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_storeTail; // @[LSQBRAM.scala 74:18:@43653.4]
  wire [3:0] GA_io_storeHead; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_storeEmpty; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_bbStart; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_bbStartSignals_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_bbStartSignals_1; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_readyToPrevious_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_readyToPrevious_1; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  GA_io_storePortsEnable_0; // @[LSQBRAM.scala 74:18:@43653.4]
  wire  LOAD_PORT_LSQ_A_clock; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_reset; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_addrFromPrev_ready; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_addrFromPrev_valid; // @[LSQBRAM.scala 77:11:@43656.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_addrFromPrev_bits; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_dataToNext_ready; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_dataToNext_valid; // @[LSQBRAM.scala 77:11:@43656.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_dataToNext_bits; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_loadAddrEnable; // @[LSQBRAM.scala 77:11:@43656.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_addrToLoadQueue; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid; // @[LSQBRAM.scala 77:11:@43656.4]
  wire [31:0] LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits; // @[LSQBRAM.scala 77:11:@43656.4]
  wire  STORE_DATA_PORT_LSQ_A_clock; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_DATA_PORT_LSQ_A_reset; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid; // @[LSQBRAM.scala 80:11:@43672.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_DATA_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_DATA_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 80:11:@43672.4]
  wire [31:0] STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 80:11:@43672.4]
  wire  STORE_ADDR_PORT_LSQ_A_clock; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  STORE_ADDR_PORT_LSQ_A_reset; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid; // @[LSQBRAM.scala 83:11:@43682.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_portEnable; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  STORE_ADDR_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 83:11:@43682.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 83:11:@43682.4]
  wire  storeEmpty; // @[LSQBRAM.scala 46:24:@43623.4 LSQBRAM.scala 151:14:@44021.4]
  wire  loadEmpty; // @[LSQBRAM.scala 52:23:@43629.4 LSQBRAM.scala 119:13:@43876.4]
  wire [15:0] storeTail; // @[LSQBRAM.scala 44:23:@43621.4 LSQBRAM.scala 149:13:@44019.4]
  wire [15:0] storeHead; // @[LSQBRAM.scala 45:23:@43622.4 LSQBRAM.scala 150:13:@44020.4]
  wire [15:0] loadTail; // @[LSQBRAM.scala 50:22:@43627.4 LSQBRAM.scala 117:12:@43874.4]
  wire [15:0] loadHead; // @[LSQBRAM.scala 51:22:@43628.4 LSQBRAM.scala 118:12:@43875.4]
  STORE_QUEUE_LSQ_A storeQ ( // @[LSQBRAM.scala 72:22:@43647.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(storeQ_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(storeQ_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(storeQ_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(storeQ_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(storeQ_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(storeQ_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(storeQ_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(storeQ_io_bbStoreOffsets_15),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadAddressDone_8(storeQ_io_loadAddressDone_8),
    .io_loadAddressDone_9(storeQ_io_loadAddressDone_9),
    .io_loadAddressDone_10(storeQ_io_loadAddressDone_10),
    .io_loadAddressDone_11(storeQ_io_loadAddressDone_11),
    .io_loadAddressDone_12(storeQ_io_loadAddressDone_12),
    .io_loadAddressDone_13(storeQ_io_loadAddressDone_13),
    .io_loadAddressDone_14(storeQ_io_loadAddressDone_14),
    .io_loadAddressDone_15(storeQ_io_loadAddressDone_15),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadDataDone_8(storeQ_io_loadDataDone_8),
    .io_loadDataDone_9(storeQ_io_loadDataDone_9),
    .io_loadDataDone_10(storeQ_io_loadDataDone_10),
    .io_loadDataDone_11(storeQ_io_loadDataDone_11),
    .io_loadDataDone_12(storeQ_io_loadDataDone_12),
    .io_loadDataDone_13(storeQ_io_loadDataDone_13),
    .io_loadDataDone_14(storeQ_io_loadDataDone_14),
    .io_loadDataDone_15(storeQ_io_loadDataDone_15),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_loadAddressQueue_8(storeQ_io_loadAddressQueue_8),
    .io_loadAddressQueue_9(storeQ_io_loadAddressQueue_9),
    .io_loadAddressQueue_10(storeQ_io_loadAddressQueue_10),
    .io_loadAddressQueue_11(storeQ_io_loadAddressQueue_11),
    .io_loadAddressQueue_12(storeQ_io_loadAddressQueue_12),
    .io_loadAddressQueue_13(storeQ_io_loadAddressQueue_13),
    .io_loadAddressQueue_14(storeQ_io_loadAddressQueue_14),
    .io_loadAddressQueue_15(storeQ_io_loadAddressQueue_15),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(storeQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(storeQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(storeQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(storeQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(storeQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(storeQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(storeQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(storeQ_io_storeAddrDone_15),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeDataDone_8(storeQ_io_storeDataDone_8),
    .io_storeDataDone_9(storeQ_io_storeDataDone_9),
    .io_storeDataDone_10(storeQ_io_storeDataDone_10),
    .io_storeDataDone_11(storeQ_io_storeDataDone_11),
    .io_storeDataDone_12(storeQ_io_storeDataDone_12),
    .io_storeDataDone_13(storeQ_io_storeDataDone_13),
    .io_storeDataDone_14(storeQ_io_storeDataDone_14),
    .io_storeDataDone_15(storeQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(storeQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(storeQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(storeQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(storeQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(storeQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(storeQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(storeQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(storeQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(storeQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(storeQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(storeQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(storeQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(storeQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(storeQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(storeQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(storeQ_io_storeDataQueue_15),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeEnableToMem(storeQ_io_storeEnableToMem),
    .io_memIsReadyForStores(storeQ_io_memIsReadyForStores)
  );
  LOAD_QUEUE_LSQ_A loadQ ( // @[LSQBRAM.scala 73:21:@43650.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(loadQ_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(loadQ_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(loadQ_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(loadQ_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(loadQ_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(loadQ_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(loadQ_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(loadQ_io_bbLoadOffsets_15),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(loadQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(loadQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(loadQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(loadQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(loadQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(loadQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(loadQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(loadQ_io_storeAddrDone_15),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeDataDone_8(loadQ_io_storeDataDone_8),
    .io_storeDataDone_9(loadQ_io_storeDataDone_9),
    .io_storeDataDone_10(loadQ_io_storeDataDone_10),
    .io_storeDataDone_11(loadQ_io_storeDataDone_11),
    .io_storeDataDone_12(loadQ_io_storeDataDone_12),
    .io_storeDataDone_13(loadQ_io_storeDataDone_13),
    .io_storeDataDone_14(loadQ_io_storeDataDone_14),
    .io_storeDataDone_15(loadQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(loadQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(loadQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(loadQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(loadQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(loadQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(loadQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(loadQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(loadQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(loadQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(loadQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(loadQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(loadQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(loadQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(loadQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(loadQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(loadQ_io_storeDataQueue_15),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadAddrDone_8(loadQ_io_loadAddrDone_8),
    .io_loadAddrDone_9(loadQ_io_loadAddrDone_9),
    .io_loadAddrDone_10(loadQ_io_loadAddrDone_10),
    .io_loadAddrDone_11(loadQ_io_loadAddrDone_11),
    .io_loadAddrDone_12(loadQ_io_loadAddrDone_12),
    .io_loadAddrDone_13(loadQ_io_loadAddrDone_13),
    .io_loadAddrDone_14(loadQ_io_loadAddrDone_14),
    .io_loadAddrDone_15(loadQ_io_loadAddrDone_15),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadDataDone_8(loadQ_io_loadDataDone_8),
    .io_loadDataDone_9(loadQ_io_loadDataDone_9),
    .io_loadDataDone_10(loadQ_io_loadDataDone_10),
    .io_loadDataDone_11(loadQ_io_loadDataDone_11),
    .io_loadDataDone_12(loadQ_io_loadDataDone_12),
    .io_loadDataDone_13(loadQ_io_loadDataDone_13),
    .io_loadDataDone_14(loadQ_io_loadDataDone_14),
    .io_loadDataDone_15(loadQ_io_loadDataDone_15),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrQueue_8(loadQ_io_loadAddrQueue_8),
    .io_loadAddrQueue_9(loadQ_io_loadAddrQueue_9),
    .io_loadAddrQueue_10(loadQ_io_loadAddrQueue_10),
    .io_loadAddrQueue_11(loadQ_io_loadAddrQueue_11),
    .io_loadAddrQueue_12(loadQ_io_loadAddrQueue_12),
    .io_loadAddrQueue_13(loadQ_io_loadAddrQueue_13),
    .io_loadAddrQueue_14(loadQ_io_loadAddrQueue_14),
    .io_loadAddrQueue_15(loadQ_io_loadAddrQueue_15),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadEnableToMem(loadQ_io_loadEnableToMem),
    .io_memIsReadyForLoads(loadQ_io_memIsReadyForLoads)
  );
  GROUP_ALLOCATOR_LSQ_A GA ( // @[LSQBRAM.scala 74:18:@43653.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(GA_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(GA_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(GA_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(GA_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(GA_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(GA_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(GA_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(GA_io_bbLoadOffsets_15),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(GA_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(GA_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(GA_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(GA_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(GA_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(GA_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(GA_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(GA_io_bbStoreOffsets_15),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_bbStartSignals_1(GA_io_bbStartSignals_1),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_readyToPrevious_1(GA_io_readyToPrevious_1),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0)
  );
  LOAD_PORT_LSQ_A LOAD_PORT_LSQ_A ( // @[LSQBRAM.scala 77:11:@43656.4]
    .clock(LOAD_PORT_LSQ_A_clock),
    .reset(LOAD_PORT_LSQ_A_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_A_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_A_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_A_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_A_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_A_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_A_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_A_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_A_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_A_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_A STORE_DATA_PORT_LSQ_A ( // @[LSQBRAM.scala 80:11:@43672.4]
    .clock(STORE_DATA_PORT_LSQ_A_clock),
    .reset(STORE_DATA_PORT_LSQ_A_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_A_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_A_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_A STORE_ADDR_PORT_LSQ_A ( // @[LSQBRAM.scala 83:11:@43682.4]
    .clock(STORE_ADDR_PORT_LSQ_A_clock),
    .reset(STORE_ADDR_PORT_LSQ_A_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_A_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_A_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 46:24:@43623.4 LSQBRAM.scala 151:14:@44021.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 52:23:@43629.4 LSQBRAM.scala 119:13:@43876.4]
  assign storeTail = {{12'd0}, storeQ_io_storeTail}; // @[LSQBRAM.scala 44:23:@43621.4 LSQBRAM.scala 149:13:@44019.4]
  assign storeHead = {{12'd0}, storeQ_io_storeHead}; // @[LSQBRAM.scala 45:23:@43622.4 LSQBRAM.scala 150:13:@44020.4]
  assign loadTail = {{12'd0}, loadQ_io_loadTail}; // @[LSQBRAM.scala 50:22:@43627.4 LSQBRAM.scala 117:12:@43874.4]
  assign loadHead = {{12'd0}, loadQ_io_loadHead}; // @[LSQBRAM.scala 51:22:@43628.4 LSQBRAM.scala 118:12:@43875.4]
  assign io_storeDataOut = storeQ_io_storeDataToMem; // @[LSQBRAM.scala 161:19:@44091.4]
  assign io_storeAddrOut = storeQ_io_storeAddrToMem; // @[LSQBRAM.scala 160:19:@44090.4]
  assign io_storeEnable = storeQ_io_storeEnableToMem; // @[LSQBRAM.scala 162:18:@44092.4]
  assign io_loadAddrOut = loadQ_io_loadAddrToMem; // @[LSQBRAM.scala 135:18:@43932.4]
  assign io_loadEnable = loadQ_io_loadEnableToMem; // @[LSQBRAM.scala 136:17:@43933.4]
  assign io_bbReadyToPrevs_0 = GA_io_readyToPrevious_0; // @[LSQBRAM.scala 102:21:@43769.4]
  assign io_bbReadyToPrevs_1 = GA_io_readyToPrevious_1; // @[LSQBRAM.scala 102:21:@43770.4]
  assign io_rdPortsPrev_0_ready = LOAD_PORT_LSQ_A_io_addrFromPrev_ready; // @[LSQBRAM.scala 166:31:@44096.4]
  assign io_rdPortsNext_0_valid = LOAD_PORT_LSQ_A_io_dataToNext_valid; // @[LSQBRAM.scala 168:23:@44099.4]
  assign io_rdPortsNext_0_bits = LOAD_PORT_LSQ_A_io_dataToNext_bits; // @[LSQBRAM.scala 168:23:@44098.4]
  assign io_wrAddrPorts_0_ready = STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 182:39:@44114.4]
  assign io_wrDataPorts_0_ready = STORE_DATA_PORT_LSQ_A_io_dataFromPrev_ready; // @[LSQBRAM.scala 177:36:@44108.4]
  assign io_Empty_Valid = storeEmpty & loadEmpty; // @[LSQBRAM.scala 86:18:@43693.4]
  assign storeQ_clock = clock; // @[:@43648.4]
  assign storeQ_reset = reset; // @[:@43649.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 145:21:@43985.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQBRAM.scala 146:28:@43986.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQBRAM.scala 146:28:@43987.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQBRAM.scala 146:28:@43988.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQBRAM.scala 146:28:@43989.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQBRAM.scala 146:28:@43990.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQBRAM.scala 146:28:@43991.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQBRAM.scala 146:28:@43992.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQBRAM.scala 146:28:@43993.4]
  assign storeQ_io_bbStoreOffsets_8 = GA_io_bbStoreOffsets_8; // @[LSQBRAM.scala 146:28:@43994.4]
  assign storeQ_io_bbStoreOffsets_9 = GA_io_bbStoreOffsets_9; // @[LSQBRAM.scala 146:28:@43995.4]
  assign storeQ_io_bbStoreOffsets_10 = GA_io_bbStoreOffsets_10; // @[LSQBRAM.scala 146:28:@43996.4]
  assign storeQ_io_bbStoreOffsets_11 = GA_io_bbStoreOffsets_11; // @[LSQBRAM.scala 146:28:@43997.4]
  assign storeQ_io_bbStoreOffsets_12 = GA_io_bbStoreOffsets_12; // @[LSQBRAM.scala 146:28:@43998.4]
  assign storeQ_io_bbStoreOffsets_13 = GA_io_bbStoreOffsets_13; // @[LSQBRAM.scala 146:28:@43999.4]
  assign storeQ_io_bbStoreOffsets_14 = GA_io_bbStoreOffsets_14; // @[LSQBRAM.scala 146:28:@44000.4]
  assign storeQ_io_bbStoreOffsets_15 = GA_io_bbStoreOffsets_15; // @[LSQBRAM.scala 146:28:@44001.4]
  assign storeQ_io_bbNumStores = GA_io_bbNumStores; // @[LSQBRAM.scala 148:25:@44018.4]
  assign storeQ_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 139:22:@43934.4]
  assign storeQ_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 140:22:@43935.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 141:23:@43936.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQBRAM.scala 142:29:@43937.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQBRAM.scala 142:29:@43938.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQBRAM.scala 142:29:@43939.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQBRAM.scala 142:29:@43940.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQBRAM.scala 142:29:@43941.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQBRAM.scala 142:29:@43942.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQBRAM.scala 142:29:@43943.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQBRAM.scala 142:29:@43944.4]
  assign storeQ_io_loadAddressDone_8 = loadQ_io_loadAddrDone_8; // @[LSQBRAM.scala 142:29:@43945.4]
  assign storeQ_io_loadAddressDone_9 = loadQ_io_loadAddrDone_9; // @[LSQBRAM.scala 142:29:@43946.4]
  assign storeQ_io_loadAddressDone_10 = loadQ_io_loadAddrDone_10; // @[LSQBRAM.scala 142:29:@43947.4]
  assign storeQ_io_loadAddressDone_11 = loadQ_io_loadAddrDone_11; // @[LSQBRAM.scala 142:29:@43948.4]
  assign storeQ_io_loadAddressDone_12 = loadQ_io_loadAddrDone_12; // @[LSQBRAM.scala 142:29:@43949.4]
  assign storeQ_io_loadAddressDone_13 = loadQ_io_loadAddrDone_13; // @[LSQBRAM.scala 142:29:@43950.4]
  assign storeQ_io_loadAddressDone_14 = loadQ_io_loadAddrDone_14; // @[LSQBRAM.scala 142:29:@43951.4]
  assign storeQ_io_loadAddressDone_15 = loadQ_io_loadAddrDone_15; // @[LSQBRAM.scala 142:29:@43952.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQBRAM.scala 143:26:@43953.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQBRAM.scala 143:26:@43954.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQBRAM.scala 143:26:@43955.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQBRAM.scala 143:26:@43956.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQBRAM.scala 143:26:@43957.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQBRAM.scala 143:26:@43958.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQBRAM.scala 143:26:@43959.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQBRAM.scala 143:26:@43960.4]
  assign storeQ_io_loadDataDone_8 = loadQ_io_loadDataDone_8; // @[LSQBRAM.scala 143:26:@43961.4]
  assign storeQ_io_loadDataDone_9 = loadQ_io_loadDataDone_9; // @[LSQBRAM.scala 143:26:@43962.4]
  assign storeQ_io_loadDataDone_10 = loadQ_io_loadDataDone_10; // @[LSQBRAM.scala 143:26:@43963.4]
  assign storeQ_io_loadDataDone_11 = loadQ_io_loadDataDone_11; // @[LSQBRAM.scala 143:26:@43964.4]
  assign storeQ_io_loadDataDone_12 = loadQ_io_loadDataDone_12; // @[LSQBRAM.scala 143:26:@43965.4]
  assign storeQ_io_loadDataDone_13 = loadQ_io_loadDataDone_13; // @[LSQBRAM.scala 143:26:@43966.4]
  assign storeQ_io_loadDataDone_14 = loadQ_io_loadDataDone_14; // @[LSQBRAM.scala 143:26:@43967.4]
  assign storeQ_io_loadDataDone_15 = loadQ_io_loadDataDone_15; // @[LSQBRAM.scala 143:26:@43968.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQBRAM.scala 144:30:@43969.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQBRAM.scala 144:30:@43970.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQBRAM.scala 144:30:@43971.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQBRAM.scala 144:30:@43972.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQBRAM.scala 144:30:@43973.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQBRAM.scala 144:30:@43974.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQBRAM.scala 144:30:@43975.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQBRAM.scala 144:30:@43976.4]
  assign storeQ_io_loadAddressQueue_8 = loadQ_io_loadAddrQueue_8; // @[LSQBRAM.scala 144:30:@43977.4]
  assign storeQ_io_loadAddressQueue_9 = loadQ_io_loadAddrQueue_9; // @[LSQBRAM.scala 144:30:@43978.4]
  assign storeQ_io_loadAddressQueue_10 = loadQ_io_loadAddrQueue_10; // @[LSQBRAM.scala 144:30:@43979.4]
  assign storeQ_io_loadAddressQueue_11 = loadQ_io_loadAddrQueue_11; // @[LSQBRAM.scala 144:30:@43980.4]
  assign storeQ_io_loadAddressQueue_12 = loadQ_io_loadAddrQueue_12; // @[LSQBRAM.scala 144:30:@43981.4]
  assign storeQ_io_loadAddressQueue_13 = loadQ_io_loadAddrQueue_13; // @[LSQBRAM.scala 144:30:@43982.4]
  assign storeQ_io_loadAddressQueue_14 = loadQ_io_loadAddrQueue_14; // @[LSQBRAM.scala 144:30:@43983.4]
  assign storeQ_io_loadAddressQueue_15 = loadQ_io_loadAddrQueue_15; // @[LSQBRAM.scala 144:30:@43984.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 156:29:@44086.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 157:32:@44087.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_A_io_storeDataEnable; // @[LSQBRAM.scala 158:29:@44088.4]
  assign storeQ_io_addressFromStorePorts_0 = STORE_ADDR_PORT_LSQ_A_io_dataToStoreQueue; // @[LSQBRAM.scala 159:35:@44089.4]
  assign storeQ_io_memIsReadyForStores = io_memIsReadyForStores; // @[LSQBRAM.scala 163:33:@44093.4]
  assign loadQ_clock = clock; // @[:@43651.4]
  assign loadQ_reset = reset; // @[:@43652.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQBRAM.scala 113:20:@43840.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQBRAM.scala 114:26:@43841.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQBRAM.scala 114:26:@43842.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQBRAM.scala 114:26:@43843.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQBRAM.scala 114:26:@43844.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQBRAM.scala 114:26:@43845.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQBRAM.scala 114:26:@43846.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQBRAM.scala 114:26:@43847.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQBRAM.scala 114:26:@43848.4]
  assign loadQ_io_bbLoadOffsets_8 = GA_io_bbLoadOffsets_8; // @[LSQBRAM.scala 114:26:@43849.4]
  assign loadQ_io_bbLoadOffsets_9 = GA_io_bbLoadOffsets_9; // @[LSQBRAM.scala 114:26:@43850.4]
  assign loadQ_io_bbLoadOffsets_10 = GA_io_bbLoadOffsets_10; // @[LSQBRAM.scala 114:26:@43851.4]
  assign loadQ_io_bbLoadOffsets_11 = GA_io_bbLoadOffsets_11; // @[LSQBRAM.scala 114:26:@43852.4]
  assign loadQ_io_bbLoadOffsets_12 = GA_io_bbLoadOffsets_12; // @[LSQBRAM.scala 114:26:@43853.4]
  assign loadQ_io_bbLoadOffsets_13 = GA_io_bbLoadOffsets_13; // @[LSQBRAM.scala 114:26:@43854.4]
  assign loadQ_io_bbLoadOffsets_14 = GA_io_bbLoadOffsets_14; // @[LSQBRAM.scala 114:26:@43855.4]
  assign loadQ_io_bbLoadOffsets_15 = GA_io_bbLoadOffsets_15; // @[LSQBRAM.scala 114:26:@43856.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQBRAM.scala 116:23:@43873.4]
  assign loadQ_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 106:22:@43773.4]
  assign loadQ_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 107:22:@43774.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 108:23:@43775.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQBRAM.scala 109:26:@43776.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQBRAM.scala 109:26:@43777.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQBRAM.scala 109:26:@43778.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQBRAM.scala 109:26:@43779.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQBRAM.scala 109:26:@43780.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQBRAM.scala 109:26:@43781.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQBRAM.scala 109:26:@43782.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQBRAM.scala 109:26:@43783.4]
  assign loadQ_io_storeAddrDone_8 = storeQ_io_storeAddrDone_8; // @[LSQBRAM.scala 109:26:@43784.4]
  assign loadQ_io_storeAddrDone_9 = storeQ_io_storeAddrDone_9; // @[LSQBRAM.scala 109:26:@43785.4]
  assign loadQ_io_storeAddrDone_10 = storeQ_io_storeAddrDone_10; // @[LSQBRAM.scala 109:26:@43786.4]
  assign loadQ_io_storeAddrDone_11 = storeQ_io_storeAddrDone_11; // @[LSQBRAM.scala 109:26:@43787.4]
  assign loadQ_io_storeAddrDone_12 = storeQ_io_storeAddrDone_12; // @[LSQBRAM.scala 109:26:@43788.4]
  assign loadQ_io_storeAddrDone_13 = storeQ_io_storeAddrDone_13; // @[LSQBRAM.scala 109:26:@43789.4]
  assign loadQ_io_storeAddrDone_14 = storeQ_io_storeAddrDone_14; // @[LSQBRAM.scala 109:26:@43790.4]
  assign loadQ_io_storeAddrDone_15 = storeQ_io_storeAddrDone_15; // @[LSQBRAM.scala 109:26:@43791.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQBRAM.scala 110:26:@43792.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQBRAM.scala 110:26:@43793.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQBRAM.scala 110:26:@43794.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQBRAM.scala 110:26:@43795.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQBRAM.scala 110:26:@43796.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQBRAM.scala 110:26:@43797.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQBRAM.scala 110:26:@43798.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQBRAM.scala 110:26:@43799.4]
  assign loadQ_io_storeDataDone_8 = storeQ_io_storeDataDone_8; // @[LSQBRAM.scala 110:26:@43800.4]
  assign loadQ_io_storeDataDone_9 = storeQ_io_storeDataDone_9; // @[LSQBRAM.scala 110:26:@43801.4]
  assign loadQ_io_storeDataDone_10 = storeQ_io_storeDataDone_10; // @[LSQBRAM.scala 110:26:@43802.4]
  assign loadQ_io_storeDataDone_11 = storeQ_io_storeDataDone_11; // @[LSQBRAM.scala 110:26:@43803.4]
  assign loadQ_io_storeDataDone_12 = storeQ_io_storeDataDone_12; // @[LSQBRAM.scala 110:26:@43804.4]
  assign loadQ_io_storeDataDone_13 = storeQ_io_storeDataDone_13; // @[LSQBRAM.scala 110:26:@43805.4]
  assign loadQ_io_storeDataDone_14 = storeQ_io_storeDataDone_14; // @[LSQBRAM.scala 110:26:@43806.4]
  assign loadQ_io_storeDataDone_15 = storeQ_io_storeDataDone_15; // @[LSQBRAM.scala 110:26:@43807.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQBRAM.scala 111:27:@43808.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQBRAM.scala 111:27:@43809.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQBRAM.scala 111:27:@43810.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQBRAM.scala 111:27:@43811.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQBRAM.scala 111:27:@43812.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQBRAM.scala 111:27:@43813.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQBRAM.scala 111:27:@43814.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQBRAM.scala 111:27:@43815.4]
  assign loadQ_io_storeAddrQueue_8 = storeQ_io_storeAddrQueue_8; // @[LSQBRAM.scala 111:27:@43816.4]
  assign loadQ_io_storeAddrQueue_9 = storeQ_io_storeAddrQueue_9; // @[LSQBRAM.scala 111:27:@43817.4]
  assign loadQ_io_storeAddrQueue_10 = storeQ_io_storeAddrQueue_10; // @[LSQBRAM.scala 111:27:@43818.4]
  assign loadQ_io_storeAddrQueue_11 = storeQ_io_storeAddrQueue_11; // @[LSQBRAM.scala 111:27:@43819.4]
  assign loadQ_io_storeAddrQueue_12 = storeQ_io_storeAddrQueue_12; // @[LSQBRAM.scala 111:27:@43820.4]
  assign loadQ_io_storeAddrQueue_13 = storeQ_io_storeAddrQueue_13; // @[LSQBRAM.scala 111:27:@43821.4]
  assign loadQ_io_storeAddrQueue_14 = storeQ_io_storeAddrQueue_14; // @[LSQBRAM.scala 111:27:@43822.4]
  assign loadQ_io_storeAddrQueue_15 = storeQ_io_storeAddrQueue_15; // @[LSQBRAM.scala 111:27:@43823.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQBRAM.scala 112:27:@43824.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQBRAM.scala 112:27:@43825.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQBRAM.scala 112:27:@43826.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQBRAM.scala 112:27:@43827.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQBRAM.scala 112:27:@43828.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQBRAM.scala 112:27:@43829.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQBRAM.scala 112:27:@43830.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQBRAM.scala 112:27:@43831.4]
  assign loadQ_io_storeDataQueue_8 = storeQ_io_storeDataQueue_8; // @[LSQBRAM.scala 112:27:@43832.4]
  assign loadQ_io_storeDataQueue_9 = storeQ_io_storeDataQueue_9; // @[LSQBRAM.scala 112:27:@43833.4]
  assign loadQ_io_storeDataQueue_10 = storeQ_io_storeDataQueue_10; // @[LSQBRAM.scala 112:27:@43834.4]
  assign loadQ_io_storeDataQueue_11 = storeQ_io_storeDataQueue_11; // @[LSQBRAM.scala 112:27:@43835.4]
  assign loadQ_io_storeDataQueue_12 = storeQ_io_storeDataQueue_12; // @[LSQBRAM.scala 112:27:@43836.4]
  assign loadQ_io_storeDataQueue_13 = storeQ_io_storeDataQueue_13; // @[LSQBRAM.scala 112:27:@43837.4]
  assign loadQ_io_storeDataQueue_14 = storeQ_io_storeDataQueue_14; // @[LSQBRAM.scala 112:27:@43838.4]
  assign loadQ_io_storeDataQueue_15 = storeQ_io_storeDataQueue_15; // @[LSQBRAM.scala 112:27:@43839.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_A_io_loadAddrEnable; // @[LSQBRAM.scala 130:32:@43929.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_A_io_addrToLoadQueue; // @[LSQBRAM.scala 129:35:@43928.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_A_io_dataFromLoadQueue_ready; // @[LSQBRAM.scala 127:33:@43927.4]
  assign loadQ_io_loadDataFromMem = io_loadDataIn; // @[LSQBRAM.scala 133:28:@43930.4]
  assign loadQ_io_memIsReadyForLoads = io_memIsReadyForLoads; // @[LSQBRAM.scala 134:31:@43931.4]
  assign GA_io_loadTail = loadTail[3:0]; // @[LSQBRAM.scala 91:18:@43727.4]
  assign GA_io_loadHead = loadHead[3:0]; // @[LSQBRAM.scala 92:18:@43728.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQBRAM.scala 93:19:@43729.4]
  assign GA_io_storeTail = storeTail[3:0]; // @[LSQBRAM.scala 97:19:@43763.4]
  assign GA_io_storeHead = storeHead[3:0]; // @[LSQBRAM.scala 98:19:@43764.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQBRAM.scala 99:20:@43765.4]
  assign GA_io_bbStartSignals_0 = io_bbpValids_0; // @[LSQBRAM.scala 101:24:@43767.4]
  assign GA_io_bbStartSignals_1 = io_bbpValids_1; // @[LSQBRAM.scala 101:24:@43768.4]
  assign LOAD_PORT_LSQ_A_clock = clock; // @[:@43657.4]
  assign LOAD_PORT_LSQ_A_reset = reset; // @[:@43658.4]
  assign LOAD_PORT_LSQ_A_io_addrFromPrev_valid = io_rdPortsPrev_0_valid; // @[LSQBRAM.scala 76:26:@43670.4]
  assign LOAD_PORT_LSQ_A_io_addrFromPrev_bits = io_rdPortsPrev_0_bits; // @[LSQBRAM.scala 76:26:@43669.4]
  assign LOAD_PORT_LSQ_A_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQBRAM.scala 76:26:@43668.4]
  assign LOAD_PORT_LSQ_A_io_dataToNext_ready = io_rdPortsNext_0_ready; // @[LSQBRAM.scala 76:26:@43667.4]
  assign LOAD_PORT_LSQ_A_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQBRAM.scala 76:26:@43661.4]
  assign LOAD_PORT_LSQ_A_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQBRAM.scala 76:26:@43660.4]
  assign STORE_DATA_PORT_LSQ_A_clock = clock; // @[:@43673.4]
  assign STORE_DATA_PORT_LSQ_A_reset = reset; // @[:@43674.4]
  assign STORE_DATA_PORT_LSQ_A_io_dataFromPrev_valid = io_wrDataPorts_0_valid; // @[LSQBRAM.scala 79:31:@43680.4]
  assign STORE_DATA_PORT_LSQ_A_io_dataFromPrev_bits = io_wrDataPorts_0_bits; // @[LSQBRAM.scala 79:31:@43679.4]
  assign STORE_DATA_PORT_LSQ_A_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 79:31:@43678.4]
  assign STORE_ADDR_PORT_LSQ_A_clock = clock; // @[:@43683.4]
  assign STORE_ADDR_PORT_LSQ_A_reset = reset; // @[:@43684.4]
  assign STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_valid = io_wrAddrPorts_0_valid; // @[LSQBRAM.scala 82:34:@43690.4]
  assign STORE_ADDR_PORT_LSQ_A_io_dataFromPrev_bits = io_wrAddrPorts_0_bits; // @[LSQBRAM.scala 82:34:@43689.4]
  assign STORE_ADDR_PORT_LSQ_A_io_portEnable = GA_io_storePortsEnable_0; // @[LSQBRAM.scala 82:34:@43688.4]
endmodule
